VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO register_file
  CLASS BLOCK ;
  FOREIGN register_file ;
  ORIGIN 0.000 0.000 ;
  SIZE 96.345 BY 107.065 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 18.655 10.640 20.255 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.930 10.640 41.530 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 61.205 10.640 62.805 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 82.480 10.640 84.080 95.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 23.920 90.860 25.520 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 45.000 90.860 46.600 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 66.080 90.860 67.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 87.160 90.860 88.760 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 15.355 10.640 16.955 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 36.630 10.640 38.230 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 57.905 10.640 59.505 95.440 ;
    END
    PORT
      LAYER met4 ;
        RECT 79.180 10.640 80.780 95.440 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 20.620 90.860 22.220 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 41.700 90.860 43.300 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 62.780 90.860 64.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 83.860 90.860 85.460 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END clk
  PIN readData1[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END readData1[0]
  PIN readData1[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END readData1[1]
  PIN readData1[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END readData1[2]
  PIN readData1[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 48.390 103.065 48.670 107.065 ;
    END
  END readData1[3]
  PIN readData1[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.345 78.240 96.345 78.840 ;
    END
  END readData1[4]
  PIN readData1[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 103.065 64.770 107.065 ;
    END
  END readData1[5]
  PIN readData1[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.345 27.240 96.345 27.840 ;
    END
  END readData1[6]
  PIN readData1[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 58.050 0.000 58.330 4.000 ;
    END
  END readData1[7]
  PIN readData2[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END readData2[0]
  PIN readData2[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END readData2[1]
  PIN readData2[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END readData2[2]
  PIN readData2[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 51.610 103.065 51.890 107.065 ;
    END
  END readData2[3]
  PIN readData2[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.345 74.840 96.345 75.440 ;
    END
  END readData2[4]
  PIN readData2[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.345 71.440 96.345 72.040 ;
    END
  END readData2[5]
  PIN readData2[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 92.345 23.840 96.345 24.440 ;
    END
  END readData2[6]
  PIN readData2[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END readData2[7]
  PIN readReg1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 92.345 30.640 96.345 31.240 ;
    END
  END readReg1[0]
  PIN readReg1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 92.345 37.440 96.345 38.040 ;
    END
  END readReg1[1]
  PIN readReg1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END readReg1[2]
  PIN readReg2[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met3 ;
        RECT 92.345 34.040 96.345 34.640 ;
    END
  END readReg2[0]
  PIN readReg2[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 92.345 40.840 96.345 41.440 ;
    END
  END readReg2[1]
  PIN readReg2[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 61.240 4.000 61.840 ;
    END
  END readReg2[2]
  PIN regWrite
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END regWrite
  PIN writeData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END writeData[0]
  PIN writeData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END writeData[1]
  PIN writeData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END writeData[2]
  PIN writeData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 45.170 103.065 45.450 107.065 ;
    END
  END writeData[3]
  PIN writeData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 92.345 64.640 96.345 65.240 ;
    END
  END writeData[4]
  PIN writeData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 92.345 51.040 96.345 51.640 ;
    END
  END writeData[5]
  PIN writeData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 92.345 17.040 96.345 17.640 ;
    END
  END writeData[6]
  PIN writeData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END writeData[7]
  PIN writeReg[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END writeReg[0]
  PIN writeReg[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 51.610 0.000 51.890 4.000 ;
    END
  END writeReg[1]
  PIN writeReg[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END writeReg[2]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 90.810 95.390 ;
      LAYER li1 ;
        RECT 5.520 10.795 90.620 95.285 ;
      LAYER met1 ;
        RECT 4.210 10.640 90.620 95.440 ;
      LAYER met2 ;
        RECT 4.230 102.785 44.890 103.770 ;
        RECT 45.730 102.785 48.110 103.770 ;
        RECT 48.950 102.785 51.330 103.770 ;
        RECT 52.170 102.785 64.210 103.770 ;
        RECT 65.050 102.785 89.150 103.770 ;
        RECT 4.230 4.280 89.150 102.785 ;
        RECT 4.230 4.000 19.130 4.280 ;
        RECT 19.970 4.000 32.010 4.280 ;
        RECT 32.850 4.000 35.230 4.280 ;
        RECT 36.070 4.000 41.670 4.280 ;
        RECT 42.510 4.000 44.890 4.280 ;
        RECT 45.730 4.000 48.110 4.280 ;
        RECT 48.950 4.000 51.330 4.280 ;
        RECT 52.170 4.000 54.550 4.280 ;
        RECT 55.390 4.000 57.770 4.280 ;
        RECT 58.610 4.000 60.990 4.280 ;
        RECT 61.830 4.000 89.150 4.280 ;
      LAYER met3 ;
        RECT 3.990 89.440 92.345 95.365 ;
        RECT 4.400 88.040 92.345 89.440 ;
        RECT 3.990 82.640 92.345 88.040 ;
        RECT 4.400 81.240 92.345 82.640 ;
        RECT 3.990 79.240 92.345 81.240 ;
        RECT 3.990 77.840 91.945 79.240 ;
        RECT 3.990 75.840 92.345 77.840 ;
        RECT 4.400 74.440 91.945 75.840 ;
        RECT 3.990 72.440 92.345 74.440 ;
        RECT 4.400 71.040 91.945 72.440 ;
        RECT 3.990 65.640 92.345 71.040 ;
        RECT 4.400 64.240 91.945 65.640 ;
        RECT 3.990 62.240 92.345 64.240 ;
        RECT 4.400 60.840 92.345 62.240 ;
        RECT 3.990 55.440 92.345 60.840 ;
        RECT 4.400 54.040 92.345 55.440 ;
        RECT 3.990 52.040 92.345 54.040 ;
        RECT 4.400 50.640 91.945 52.040 ;
        RECT 3.990 48.640 92.345 50.640 ;
        RECT 4.400 47.240 92.345 48.640 ;
        RECT 3.990 41.840 92.345 47.240 ;
        RECT 3.990 40.440 91.945 41.840 ;
        RECT 3.990 38.440 92.345 40.440 ;
        RECT 3.990 37.040 91.945 38.440 ;
        RECT 3.990 35.040 92.345 37.040 ;
        RECT 3.990 33.640 91.945 35.040 ;
        RECT 3.990 31.640 92.345 33.640 ;
        RECT 3.990 30.240 91.945 31.640 ;
        RECT 3.990 28.240 92.345 30.240 ;
        RECT 3.990 26.840 91.945 28.240 ;
        RECT 3.990 24.840 92.345 26.840 ;
        RECT 3.990 23.440 91.945 24.840 ;
        RECT 3.990 18.040 92.345 23.440 ;
        RECT 3.990 16.640 91.945 18.040 ;
        RECT 3.990 10.715 92.345 16.640 ;
      LAYER met4 ;
        RECT 17.775 28.735 18.255 88.905 ;
        RECT 20.655 28.735 36.230 88.905 ;
        RECT 38.630 28.735 39.530 88.905 ;
        RECT 41.930 28.735 57.505 88.905 ;
        RECT 59.905 28.735 60.805 88.905 ;
        RECT 63.205 28.735 72.385 88.905 ;
  END
END register_file
END LIBRARY

