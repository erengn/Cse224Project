* NGSPICE file created from register_file.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt register_file VGND VPWR clk readData1[0] readData1[1] readData1[2] readData1[3]
+ readData1[4] readData1[5] readData1[6] readData1[7] readData2[0] readData2[1] readData2[2]
+ readData2[3] readData2[4] readData2[5] readData2[6] readData2[7] readReg1[0] readReg1[1]
+ readReg1[2] readReg2[0] readReg2[1] readReg2[2] regWrite writeData[0] writeData[1]
+ writeData[2] writeData[3] writeData[4] writeData[5] writeData[6] writeData[7] writeReg[0]
+ writeReg[1] writeReg[2]
XTAP_TAPCELL_ROW_24_139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_501_ clknet_3_3__leaf_clk _019_ VGND VGND VPWR VPWR registers\[4\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_432_ _206_ VGND VGND VPWR VPWR _040_ sky130_fd_sc_hd__clkbuf_1
X_294_ registers\[0\]\[0\] _116_ _112_ VGND VGND VPWR VPWR _117_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_363_ net35 net9 _167_ VGND VGND VPWR VPWR _169_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_19_Left_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_415_ net43 net9 _195_ VGND VGND VPWR VPWR _197_ sky130_fd_sc_hd__mux2_1
X_346_ _159_ VGND VGND VPWR VPWR _001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_277_ _072_ registers\[0\]\[6\] net5 VGND VGND VPWR VPWR _102_ sky130_fd_sc_hd__o21ba_1
XPHY_EDGE_ROW_4_Left_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_329_ registers\[4\]\[6\] registers\[5\]\[6\] registers\[6\]\[6\] registers\[7\]\[6\]
+ _111_ _112_ VGND VGND VPWR VPWR _146_ sky130_fd_sc_hd__mux4_1
XFILLER_0_10_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold63 registers\[0\]\[3\] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 registers\[4\]\[1\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 registers\[4\]\[7\] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 registers\[3\]\[6\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_27_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput31 net31 VGND VGND VPWR VPWR readData2[4] sky130_fd_sc_hd__buf_2
Xoutput20 net20 VGND VGND VPWR VPWR readData1[1] sky130_fd_sc_hd__buf_2
XFILLER_0_27_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_362_ _168_ VGND VGND VPWR VPWR _008_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_431_ net8 net92 _205_ VGND VGND VPWR VPWR _206_ sky130_fd_sc_hd__mux2_1
X_500_ clknet_3_1__leaf_clk _018_ VGND VGND VPWR VPWR registers\[4\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_293_ net1 VGND VGND VPWR VPWR _116_ sky130_fd_sc_hd__buf_2
XFILLER_0_13_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_414_ _196_ VGND VGND VPWR VPWR _032_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_20_Left_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_345_ net73 net9 _157_ VGND VGND VPWR VPWR _159_ sky130_fd_sc_hd__mux2_1
X_276_ registers\[1\]\[6\] _070_ VGND VGND VPWR VPWR _101_ sky130_fd_sc_hd__or2b_1
XTAP_TAPCELL_ROW_8_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_328_ _110_ _141_ _145_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__o21a_1
X_259_ _070_ registers\[0\]\[3\] net5 VGND VGND VPWR VPWR _087_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold42 registers\[2\]\[6\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 registers\[7\]\[7\] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 registers\[2\]\[7\] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 registers\[6\]\[2\] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 registers\[0\]\[7\] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput32 net32 VGND VGND VPWR VPWR readData2[5] sky130_fd_sc_hd__buf_2
Xoutput21 net21 VGND VGND VPWR VPWR readData1[2] sky130_fd_sc_hd__buf_2
XFILLER_0_27_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_361_ net50 net8 _167_ VGND VGND VPWR VPWR _168_ sky130_fd_sc_hd__mux2_1
X_292_ registers\[1\]\[0\] _111_ VGND VGND VPWR VPWR _115_ sky130_fd_sc_hd__or2b_1
X_430_ _204_ VGND VGND VPWR VPWR _205_ sky130_fd_sc_hd__clkbuf_4
X_344_ _158_ VGND VGND VPWR VPWR _000_ sky130_fd_sc_hd__clkbuf_1
X_413_ net41 net8 _195_ VGND VGND VPWR VPWR _196_ sky130_fd_sc_hd__mux2_1
X_275_ registers\[4\]\[6\] registers\[5\]\[6\] registers\[6\]\[6\] registers\[7\]\[6\]
+ _065_ _066_ VGND VGND VPWR VPWR _100_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_11_100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_258_ registers\[1\]\[3\] _070_ VGND VGND VPWR VPWR _086_ sky130_fd_sc_hd__or2b_1
X_327_ _142_ _143_ _144_ _113_ net3 VGND VGND VPWR VPWR _145_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold21 registers\[2\]\[4\] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 registers\[2\]\[3\] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 registers\[3\]\[4\] VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold32 registers\[1\]\[6\] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 registers\[6\]\[7\] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput22 net22 VGND VGND VPWR VPWR readData1[3] sky130_fd_sc_hd__clkbuf_4
Xoutput33 net33 VGND VGND VPWR VPWR readData2[6] sky130_fd_sc_hd__buf_2
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_291_ registers\[4\]\[0\] registers\[5\]\[0\] registers\[6\]\[0\] registers\[7\]\[0\]
+ _111_ _113_ VGND VGND VPWR VPWR _114_ sky130_fd_sc_hd__mux4_1
X_360_ _166_ VGND VGND VPWR VPWR _167_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_489_ clknet_3_1__leaf_clk _007_ VGND VGND VPWR VPWR registers\[6\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_343_ net36 net8 _157_ VGND VGND VPWR VPWR _158_ sky130_fd_sc_hd__mux2_1
X_274_ _064_ _095_ _099_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__o21a_1
X_412_ net18 net16 net7 net17 VGND VGND VPWR VPWR _195_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_257_ registers\[4\]\[3\] registers\[5\]\[3\] registers\[6\]\[3\] registers\[7\]\[3\]
+ _065_ _066_ VGND VGND VPWR VPWR _085_ sky130_fd_sc_hd__mux4_1
X_326_ registers\[2\]\[5\] registers\[3\]\[5\] _118_ VGND VGND VPWR VPWR _144_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_8_Left_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_309_ _127_ _128_ _129_ _113_ net3 VGND VGND VPWR VPWR _130_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold11 registers\[5\]\[5\] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 registers\[7\]\[3\] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 registers\[1\]\[0\] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 registers\[4\]\[2\] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 registers\[1\]\[2\] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlygate4sd3_1
Xoutput23 net23 VGND VGND VPWR VPWR readData1[4] sky130_fd_sc_hd__buf_2
Xoutput34 net34 VGND VGND VPWR VPWR readData2[7] sky130_fd_sc_hd__buf_2
XFILLER_0_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_290_ _112_ VGND VGND VPWR VPWR _113_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_488_ clknet_3_4__leaf_clk _006_ VGND VGND VPWR VPWR registers\[6\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_273_ _096_ _097_ _098_ _067_ net6 VGND VGND VPWR VPWR _099_ sky130_fd_sc_hd__a221o_1
X_342_ _156_ VGND VGND VPWR VPWR _157_ sky130_fd_sc_hd__clkbuf_4
X_411_ _194_ VGND VGND VPWR VPWR _031_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_24_Left_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_325_ registers\[0\]\[5\] _118_ net2 VGND VGND VPWR VPWR _143_ sky130_fd_sc_hd__o21ba_1
X_256_ _064_ _080_ _084_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__o21a_1
XFILLER_0_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload0 clknet_3_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_308_ registers\[2\]\[2\] registers\[3\]\[2\] _118_ VGND VGND VPWR VPWR _129_ sky130_fd_sc_hd__mux2_1
X_239_ net4 VGND VGND VPWR VPWR _070_ sky130_fd_sc_hd__buf_2
Xhold34 registers\[4\]\[3\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 registers\[1\]\[5\] VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 registers\[3\]\[1\] VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 registers\[5\]\[2\] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 registers\[3\]\[7\] VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput24 net24 VGND VGND VPWR VPWR readData1[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_11_Left_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_487_ clknet_3_6__leaf_clk _005_ VGND VGND VPWR VPWR registers\[6\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_13_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_272_ registers\[2\]\[5\] registers\[3\]\[5\] _072_ VGND VGND VPWR VPWR _098_ sky130_fd_sc_hd__mux2_1
X_410_ net90 net15 _186_ VGND VGND VPWR VPWR _194_ sky130_fd_sc_hd__mux2_1
X_341_ net16 net7 net18 net17 VGND VGND VPWR VPWR _156_ sky130_fd_sc_hd__and4b_1
X_539_ clknet_3_0__leaf_clk _057_ VGND VGND VPWR VPWR registers\[7\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_324_ registers\[1\]\[5\] _116_ VGND VGND VPWR VPWR _142_ sky130_fd_sc_hd__or2b_1
X_255_ _081_ _082_ _083_ _067_ net6 VGND VGND VPWR VPWR _084_ sky130_fd_sc_hd__a221o_1
XFILLER_0_27_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_92 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload1 clknet_3_1__leaf_clk VGND VGND VPWR VPWR clkload1/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_21_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_238_ registers\[1\]\[0\] _065_ VGND VGND VPWR VPWR _069_ sky130_fd_sc_hd__or2b_1
X_307_ registers\[0\]\[2\] _116_ _112_ VGND VGND VPWR VPWR _128_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_30_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold46 registers\[4\]\[5\] VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 registers\[6\]\[4\] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 registers\[1\]\[3\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold57 registers\[0\]\[5\] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlygate4sd3_1
Xhold13 registers\[2\]\[2\] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput25 net25 VGND VGND VPWR VPWR readData1[6] sky130_fd_sc_hd__buf_2
XFILLER_0_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_486_ clknet_3_6__leaf_clk _004_ VGND VGND VPWR VPWR registers\[6\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_1_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_538_ clknet_3_2__leaf_clk _056_ VGND VGND VPWR VPWR registers\[7\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_271_ _072_ registers\[0\]\[5\] net5 VGND VGND VPWR VPWR _097_ sky130_fd_sc_hd__o21ba_1
X_340_ _110_ _151_ _155_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__o21a_1
X_469_ _226_ VGND VGND VPWR VPWR _057_ sky130_fd_sc_hd__clkbuf_1
X_323_ registers\[4\]\[5\] registers\[5\]\[5\] registers\[6\]\[5\] registers\[7\]\[5\]
+ _111_ _112_ VGND VGND VPWR VPWR _141_ sky130_fd_sc_hd__mux4_1
X_254_ registers\[2\]\[2\] registers\[3\]\[2\] _072_ VGND VGND VPWR VPWR _083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_9_93 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload2 clknet_3_2__leaf_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_4
X_237_ registers\[4\]\[0\] registers\[5\]\[0\] registers\[6\]\[0\] registers\[7\]\[0\]
+ _065_ _067_ VGND VGND VPWR VPWR _068_ sky130_fd_sc_hd__mux4_1
X_306_ registers\[1\]\[2\] _116_ VGND VGND VPWR VPWR _127_ sky130_fd_sc_hd__or2b_1
Xhold47 registers\[7\]\[4\] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 registers\[3\]\[0\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 registers\[0\]\[0\] VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 registers\[7\]\[2\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__dlygate4sd3_1
Xhold14 registers\[6\]\[6\] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput26 net26 VGND VGND VPWR VPWR readData1[7] sky130_fd_sc_hd__buf_2
XFILLER_0_27_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_23_135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_88 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_485_ clknet_3_3__leaf_clk _003_ VGND VGND VPWR VPWR registers\[6\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_20_127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_270_ registers\[1\]\[5\] _070_ VGND VGND VPWR VPWR _096_ sky130_fd_sc_hd__or2b_1
X_399_ _188_ VGND VGND VPWR VPWR _025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_537_ clknet_3_1__leaf_clk _055_ VGND VGND VPWR VPWR registers\[1\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_468_ net53 net9 _224_ VGND VGND VPWR VPWR _226_ sky130_fd_sc_hd__mux2_1
X_322_ _110_ _136_ _140_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__o21a_1
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_253_ _070_ registers\[0\]\[2\] _066_ VGND VGND VPWR VPWR _082_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_9_94 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload3 clknet_3_4__leaf_clk VGND VGND VPWR VPWR clkload3/Y sky130_fd_sc_hd__bufinv_16
XPHY_EDGE_ROW_28_Left_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_305_ registers\[4\]\[2\] registers\[5\]\[2\] registers\[6\]\[2\] registers\[7\]\[2\]
+ _111_ _112_ VGND VGND VPWR VPWR _126_ sky130_fd_sc_hd__mux4_1
X_236_ _066_ VGND VGND VPWR VPWR _067_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold15 registers\[7\]\[5\] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 registers\[5\]\[4\] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 registers\[7\]\[0\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 registers\[0\]\[4\] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 registers\[3\]\[2\] VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_29_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput27 net27 VGND VGND VPWR VPWR readData2[0] sky130_fd_sc_hd__buf_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_23_136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_15_Left_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_484_ clknet_3_0__leaf_clk _002_ VGND VGND VPWR VPWR registers\[6\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_467_ _225_ VGND VGND VPWR VPWR _056_ sky130_fd_sc_hd__clkbuf_1
X_398_ net79 net9 _186_ VGND VGND VPWR VPWR _188_ sky130_fd_sc_hd__mux2_1
X_536_ clknet_3_4__leaf_clk _054_ VGND VGND VPWR VPWR registers\[1\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_321_ _137_ _138_ _139_ _113_ net3 VGND VGND VPWR VPWR _140_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_0_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_252_ registers\[1\]\[2\] _070_ VGND VGND VPWR VPWR _081_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_519_ clknet_3_7__leaf_clk _037_ VGND VGND VPWR VPWR registers\[2\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_235_ net5 VGND VGND VPWR VPWR _066_ sky130_fd_sc_hd__clkbuf_4
X_304_ _110_ _121_ _125_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__o21a_1
XPHY_EDGE_ROW_3_Left_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload4 clknet_3_5__leaf_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold16 registers\[5\]\[0\] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 registers\[3\]\[5\] VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 registers\[4\]\[6\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 registers\[1\]\[7\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_95 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput28 net28 VGND VGND VPWR VPWR readData2[1] sky130_fd_sc_hd__buf_2
XFILLER_0_7_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_26_145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_483_ clknet_3_0__leaf_clk _001_ VGND VGND VPWR VPWR registers\[6\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_466_ net60 net8 _224_ VGND VGND VPWR VPWR _225_ sky130_fd_sc_hd__mux2_1
X_397_ _187_ VGND VGND VPWR VPWR _024_ sky130_fd_sc_hd__clkbuf_1
X_535_ clknet_3_6__leaf_clk _053_ VGND VGND VPWR VPWR registers\[1\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_5_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_320_ registers\[2\]\[4\] registers\[3\]\[4\] _118_ VGND VGND VPWR VPWR _139_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_251_ registers\[4\]\[2\] registers\[5\]\[2\] registers\[6\]\[2\] registers\[7\]\[2\]
+ _065_ _066_ VGND VGND VPWR VPWR _080_ sky130_fd_sc_hd__mux4_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_518_ clknet_3_7__leaf_clk _036_ VGND VGND VPWR VPWR registers\[2\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_449_ _215_ VGND VGND VPWR VPWR _048_ sky130_fd_sc_hd__clkbuf_1
Xclkload5 clknet_3_6__leaf_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_18_112 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_303_ _122_ _123_ _124_ _113_ net3 VGND VGND VPWR VPWR _125_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_234_ net4 VGND VGND VPWR VPWR _065_ sky130_fd_sc_hd__buf_4
XFILLER_0_30_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold28 registers\[5\]\[3\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 registers\[6\]\[1\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 registers\[5\]\[7\] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_10_96 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput29 net29 VGND VGND VPWR VPWR readData2[2] sky130_fd_sc_hd__buf_2
XFILLER_0_11_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_482_ clknet_3_2__leaf_clk _000_ VGND VGND VPWR VPWR registers\[6\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_3_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_534_ clknet_3_6__leaf_clk _052_ VGND VGND VPWR VPWR registers\[1\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_396_ net70 net8 _186_ VGND VGND VPWR VPWR _187_ sky130_fd_sc_hd__mux2_1
X_465_ _223_ VGND VGND VPWR VPWR _224_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_250_ _064_ _075_ _079_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__o21a_1
XFILLER_0_27_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_379_ _177_ VGND VGND VPWR VPWR _016_ sky130_fd_sc_hd__clkbuf_1
X_517_ clknet_3_3__leaf_clk _035_ VGND VGND VPWR VPWR registers\[2\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_448_ net56 net8 _214_ VGND VGND VPWR VPWR _215_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload6 clknet_3_7__leaf_clk VGND VGND VPWR VPWR clkload6/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_18_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_233_ net6 VGND VGND VPWR VPWR _064_ sky130_fd_sc_hd__inv_2
X_302_ registers\[2\]\[1\] registers\[3\]\[1\] _118_ VGND VGND VPWR VPWR _124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold29 registers\[1\]\[4\] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 registers\[2\]\[5\] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_10_97 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput19 net19 VGND VGND VPWR VPWR readData1[0] sky130_fd_sc_hd__buf_2
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_481_ _232_ VGND VGND VPWR VPWR _063_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_533_ clknet_3_3__leaf_clk _051_ VGND VGND VPWR VPWR registers\[1\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_464_ net18 net17 net16 net7 VGND VGND VPWR VPWR _223_ sky130_fd_sc_hd__and4_1
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_395_ _185_ VGND VGND VPWR VPWR _186_ sky130_fd_sc_hd__clkbuf_4
X_378_ net84 net8 _176_ VGND VGND VPWR VPWR _177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_0_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_516_ clknet_3_0__leaf_clk _034_ VGND VGND VPWR VPWR registers\[2\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_447_ net18 net17 net16 net7 VGND VGND VPWR VPWR _214_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_24_106 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_301_ registers\[0\]\[1\] _116_ _112_ VGND VGND VPWR VPWR _123_ sky130_fd_sc_hd__o21ba_1
Xhold19 registers\[7\]\[1\] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_7_Left_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_480_ net54 net15 _224_ VGND VGND VPWR VPWR _232_ sky130_fd_sc_hd__mux2_1
X_463_ _222_ VGND VGND VPWR VPWR _055_ sky130_fd_sc_hd__clkbuf_1
X_532_ clknet_3_0__leaf_clk _050_ VGND VGND VPWR VPWR registers\[1\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_394_ net18 net17 net16 net7 VGND VGND VPWR VPWR _185_ sky130_fd_sc_hd__and4b_1
XFILLER_0_14_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_515_ clknet_3_2__leaf_clk _033_ VGND VGND VPWR VPWR registers\[2\]\[1\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_446_ _213_ VGND VGND VPWR VPWR _047_ sky130_fd_sc_hd__clkbuf_1
X_377_ net17 net16 net7 net18 VGND VGND VPWR VPWR _176_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_26_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_300_ registers\[1\]\[1\] _111_ VGND VGND VPWR VPWR _122_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_23_Left_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_429_ net18 net17 net16 net7 VGND VGND VPWR VPWR _204_ sky130_fd_sc_hd__or4b_1
Xinput1 readReg1[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_2_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_10_Left_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_531_ clknet_3_2__leaf_clk _049_ VGND VGND VPWR VPWR registers\[1\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_393_ _184_ VGND VGND VPWR VPWR _023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_462_ net61 net15 _214_ VGND VGND VPWR VPWR _222_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_514_ clknet_3_2__leaf_clk _032_ VGND VGND VPWR VPWR registers\[2\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_376_ _175_ VGND VGND VPWR VPWR _015_ sky130_fd_sc_hd__clkbuf_1
X_445_ net15 net98 _205_ VGND VGND VPWR VPWR _213_ sky130_fd_sc_hd__mux2_1
X_359_ net17 net16 net7 net18 VGND VGND VPWR VPWR _166_ sky130_fd_sc_hd__and4b_1
X_428_ _203_ VGND VGND VPWR VPWR _039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput2 readReg1[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_14_109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_530_ clknet_3_2__leaf_clk _048_ VGND VGND VPWR VPWR registers\[1\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_461_ _221_ VGND VGND VPWR VPWR _054_ sky130_fd_sc_hd__clkbuf_1
X_392_ net75 net15 _176_ VGND VGND VPWR VPWR _184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_444_ _212_ VGND VGND VPWR VPWR _046_ sky130_fd_sc_hd__clkbuf_1
X_375_ net51 net15 _167_ VGND VGND VPWR VPWR _175_ sky130_fd_sc_hd__mux2_1
X_513_ clknet_3_5__leaf_clk _031_ VGND VGND VPWR VPWR registers\[3\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_358_ _165_ VGND VGND VPWR VPWR _007_ sky130_fd_sc_hd__clkbuf_1
X_427_ net87 net15 _195_ VGND VGND VPWR VPWR _203_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput3 readReg1[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_289_ net2 VGND VGND VPWR VPWR _112_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_391_ _183_ VGND VGND VPWR VPWR _022_ sky130_fd_sc_hd__clkbuf_1
X_460_ net66 net14 _214_ VGND VGND VPWR VPWR _221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_374_ _174_ VGND VGND VPWR VPWR _014_ sky130_fd_sc_hd__clkbuf_1
X_512_ clknet_3_5__leaf_clk _030_ VGND VGND VPWR VPWR registers\[3\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_443_ net14 net96 _205_ VGND VGND VPWR VPWR _212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_426_ _202_ VGND VGND VPWR VPWR _038_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_357_ net44 net15 _157_ VGND VGND VPWR VPWR _165_ sky130_fd_sc_hd__mux2_1
X_288_ net1 VGND VGND VPWR VPWR _111_ sky130_fd_sc_hd__buf_4
Xinput4 readReg2[0] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dlymetal6s2s_1
XPHY_EDGE_ROW_27_Left_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_409_ _193_ VGND VGND VPWR VPWR _030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_25_141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_14_Left_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_390_ net72 net14 _176_ VGND VGND VPWR VPWR _183_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_511_ clknet_3_7__leaf_clk _029_ VGND VGND VPWR VPWR registers\[3\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_442_ _211_ VGND VGND VPWR VPWR _045_ sky130_fd_sc_hd__clkbuf_1
X_373_ net74 net14 _167_ VGND VGND VPWR VPWR _174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_287_ net3 VGND VGND VPWR VPWR _110_ sky130_fd_sc_hd__inv_2
X_425_ net76 net14 _195_ VGND VGND VPWR VPWR _202_ sky130_fd_sc_hd__mux2_1
X_356_ _164_ VGND VGND VPWR VPWR _006_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput5 readReg2[1] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_28_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_2_Left_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_408_ net86 net14 _186_ VGND VGND VPWR VPWR _193_ sky130_fd_sc_hd__mux2_1
X_339_ _152_ _153_ _154_ _113_ net3 VGND VGND VPWR VPWR _155_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_25_142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_372_ _173_ VGND VGND VPWR VPWR _013_ sky130_fd_sc_hd__clkbuf_1
X_510_ clknet_3_7__leaf_clk _028_ VGND VGND VPWR VPWR registers\[3\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_441_ net13 net91 _205_ VGND VGND VPWR VPWR _211_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_424_ _201_ VGND VGND VPWR VPWR _037_ sky130_fd_sc_hd__clkbuf_1
X_355_ net48 net14 _157_ VGND VGND VPWR VPWR _164_ sky130_fd_sc_hd__mux2_1
X_286_ _064_ _105_ _109_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__o21a_1
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput6 readReg2[2] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_28_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_269_ registers\[4\]\[5\] registers\[5\]\[5\] registers\[6\]\[5\] registers\[7\]\[5\]
+ _065_ _066_ VGND VGND VPWR VPWR _095_ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_407_ _192_ VGND VGND VPWR VPWR _029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_338_ registers\[2\]\[7\] registers\[3\]\[7\] net1 VGND VGND VPWR VPWR _154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_371_ net45 net13 _167_ VGND VGND VPWR VPWR _173_ sky130_fd_sc_hd__mux2_1
X_440_ _210_ VGND VGND VPWR VPWR _044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_354_ _163_ VGND VGND VPWR VPWR _005_ sky130_fd_sc_hd__clkbuf_1
X_423_ net52 net13 _195_ VGND VGND VPWR VPWR _201_ sky130_fd_sc_hd__mux2_1
X_285_ _106_ _107_ _108_ _067_ net6 VGND VGND VPWR VPWR _109_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput7 regWrite VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_9_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_268_ _064_ _090_ _094_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__o21a_1
X_406_ net83 net13 _186_ VGND VGND VPWR VPWR _192_ sky130_fd_sc_hd__mux2_1
X_337_ registers\[0\]\[7\] _118_ net2 VGND VGND VPWR VPWR _153_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_11_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput10 writeData[2] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_18_Left_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_370_ _172_ VGND VGND VPWR VPWR _012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_499_ clknet_3_1__leaf_clk _017_ VGND VGND VPWR VPWR registers\[4\]\[1\] sky130_fd_sc_hd__dfxtp_1
X_353_ net42 net13 _157_ VGND VGND VPWR VPWR _163_ sky130_fd_sc_hd__mux2_1
X_422_ _200_ VGND VGND VPWR VPWR _036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_284_ registers\[2\]\[7\] registers\[3\]\[7\] net4 VGND VGND VPWR VPWR _108_ sky130_fd_sc_hd__mux2_1
Xinput8 writeData[0] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_267_ _091_ _092_ _093_ _067_ net6 VGND VGND VPWR VPWR _094_ sky130_fd_sc_hd__a221o_1
X_405_ _191_ VGND VGND VPWR VPWR _028_ sky130_fd_sc_hd__clkbuf_1
X_336_ registers\[1\]\[7\] _116_ VGND VGND VPWR VPWR _152_ sky130_fd_sc_hd__or2b_1
XFILLER_0_11_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_6_Left_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput11 writeData[3] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_2
X_319_ registers\[0\]\[4\] _118_ net2 VGND VGND VPWR VPWR _138_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_13_104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_9_Left_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_498_ clknet_3_3__leaf_clk _016_ VGND VGND VPWR VPWR registers\[4\]\[0\] sky130_fd_sc_hd__dfxtp_1
X_421_ net55 net12 _195_ VGND VGND VPWR VPWR _200_ sky130_fd_sc_hd__mux2_1
X_352_ _162_ VGND VGND VPWR VPWR _004_ sky130_fd_sc_hd__clkbuf_1
Xinput9 writeData[1] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_2
X_283_ _072_ registers\[0\]\[7\] net5 VGND VGND VPWR VPWR _107_ sky130_fd_sc_hd__o21ba_1
X_266_ registers\[2\]\[4\] registers\[3\]\[4\] _072_ VGND VGND VPWR VPWR _093_ sky130_fd_sc_hd__mux2_1
X_404_ net88 net12 _186_ VGND VGND VPWR VPWR _191_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_335_ registers\[4\]\[7\] registers\[5\]\[7\] registers\[6\]\[7\] registers\[7\]\[7\]
+ _111_ _112_ VGND VGND VPWR VPWR _151_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_22_Left_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput12 writeData[4] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
X_318_ registers\[1\]\[4\] _116_ VGND VGND VPWR VPWR _137_ sky130_fd_sc_hd__or2b_1
X_249_ _076_ _077_ _078_ _067_ net6 VGND VGND VPWR VPWR _079_ sky130_fd_sc_hd__a221o_1
XTAP_TAPCELL_ROW_16_113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_30_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_13_105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold1 registers\[5\]\[1\] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dlygate4sd3_1
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_497_ clknet_3_1__leaf_clk _015_ VGND VGND VPWR VPWR registers\[5\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_17_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_420_ _199_ VGND VGND VPWR VPWR _035_ sky130_fd_sc_hd__clkbuf_1
X_351_ net69 net12 _157_ VGND VGND VPWR VPWR _162_ sky130_fd_sc_hd__mux2_1
X_282_ registers\[1\]\[7\] _070_ VGND VGND VPWR VPWR _106_ sky130_fd_sc_hd__or2b_1
X_403_ _190_ VGND VGND VPWR VPWR _027_ sky130_fd_sc_hd__clkbuf_1
X_334_ _110_ _146_ _150_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__o21a_1
XFILLER_0_9_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_265_ _072_ registers\[0\]\[4\] net5 VGND VGND VPWR VPWR _092_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_317_ registers\[4\]\[4\] registers\[5\]\[4\] registers\[6\]\[4\] registers\[7\]\[4\]
+ _111_ _112_ VGND VGND VPWR VPWR _136_ sky130_fd_sc_hd__mux4_1
XTAP_TAPCELL_ROW_16_114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_248_ registers\[2\]\[1\] registers\[3\]\[1\] _072_ VGND VGND VPWR VPWR _078_ sky130_fd_sc_hd__mux2_1
Xinput13 writeData[5] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_7_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold2 registers\[6\]\[0\] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dlygate4sd3_1
X_496_ clknet_3_4__leaf_clk _014_ VGND VGND VPWR VPWR registers\[5\]\[6\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_350_ _161_ VGND VGND VPWR VPWR _003_ sky130_fd_sc_hd__clkbuf_1
X_281_ registers\[4\]\[7\] registers\[5\]\[7\] registers\[6\]\[7\] registers\[7\]\[7\]
+ _065_ _066_ VGND VGND VPWR VPWR _105_ sky130_fd_sc_hd__mux4_1
XFILLER_0_11_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_479_ _231_ VGND VGND VPWR VPWR _062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_402_ net85 net11 _186_ VGND VGND VPWR VPWR _190_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_264_ registers\[1\]\[4\] _070_ VGND VGND VPWR VPWR _091_ sky130_fd_sc_hd__or2b_1
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_333_ _147_ _148_ _149_ _113_ net3 VGND VGND VPWR VPWR _150_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_316_ _110_ _131_ _135_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__o21a_1
XTAP_TAPCELL_ROW_16_115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_247_ _070_ registers\[0\]\[1\] _066_ VGND VGND VPWR VPWR _077_ sky130_fd_sc_hd__o21ba_1
Xinput14 writeData[6] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_7_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold3 registers\[6\]\[3\] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_495_ clknet_3_6__leaf_clk _013_ VGND VGND VPWR VPWR registers\[5\]\[5\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_280_ _064_ _100_ _104_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__o21a_1
XFILLER_0_11_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_478_ net38 net14 _224_ VGND VGND VPWR VPWR _231_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_263_ registers\[4\]\[4\] registers\[5\]\[4\] registers\[6\]\[4\] registers\[7\]\[4\]
+ _065_ _066_ VGND VGND VPWR VPWR _090_ sky130_fd_sc_hd__mux4_1
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_401_ _189_ VGND VGND VPWR VPWR _026_ sky130_fd_sc_hd__clkbuf_1
X_332_ registers\[2\]\[6\] registers\[3\]\[6\] net1 VGND VGND VPWR VPWR _149_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_19_124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_11_98 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_26_Left_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_315_ _132_ _133_ _134_ _113_ net3 VGND VGND VPWR VPWR _135_ sky130_fd_sc_hd__a221o_1
X_246_ registers\[1\]\[1\] _065_ VGND VGND VPWR VPWR _076_ sky130_fd_sc_hd__or2b_1
Xinput15 writeData[7] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_21_130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_30_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold4 registers\[7\]\[6\] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_4_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_29_Left_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Left_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_494_ clknet_3_7__leaf_clk _012_ VGND VGND VPWR VPWR registers\[5\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_477_ _230_ VGND VGND VPWR VPWR _061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_262_ _064_ _085_ _089_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__o21a_1
X_400_ net82 net10 _186_ VGND VGND VPWR VPWR _189_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_331_ registers\[0\]\[6\] _118_ net2 VGND VGND VPWR VPWR _148_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_529_ clknet_3_4__leaf_clk _047_ VGND VGND VPWR VPWR registers\[0\]\[7\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_1_Left_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_99 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_314_ registers\[2\]\[3\] registers\[3\]\[3\] _118_ VGND VGND VPWR VPWR _134_ sky130_fd_sc_hd__mux2_1
Xinput16 writeReg[0] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dlymetal6s2s_1
X_245_ registers\[4\]\[1\] registers\[5\]\[1\] registers\[6\]\[1\] registers\[7\]\[1\]
+ _065_ _067_ VGND VGND VPWR VPWR _075_ sky130_fd_sc_hd__mux4_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold5 registers\[4\]\[4\] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_30_Left_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_493_ clknet_3_3__leaf_clk _011_ VGND VGND VPWR VPWR registers\[5\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_19_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_476_ net49 net13 _224_ VGND VGND VPWR VPWR _230_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_1_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_545_ clknet_3_1__leaf_clk _063_ VGND VGND VPWR VPWR registers\[7\]\[7\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_261_ _086_ _087_ _088_ _067_ net6 VGND VGND VPWR VPWR _089_ sky130_fd_sc_hd__a221o_1
X_330_ registers\[1\]\[6\] _116_ VGND VGND VPWR VPWR _147_ sky130_fd_sc_hd__or2b_1
X_459_ _220_ VGND VGND VPWR VPWR _053_ sky130_fd_sc_hd__clkbuf_1
X_528_ clknet_3_5__leaf_clk _046_ VGND VGND VPWR VPWR registers\[0\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_244_ _064_ _068_ _074_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__o21a_1
X_313_ registers\[0\]\[3\] _116_ net2 VGND VGND VPWR VPWR _133_ sky130_fd_sc_hd__o21ba_1
Xinput17 writeReg[1] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_2_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_84 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold6 registers\[1\]\[1\] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_492_ clknet_3_0__leaf_clk _010_ VGND VGND VPWR VPWR registers\[5\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_475_ _229_ VGND VGND VPWR VPWR _060_ sky130_fd_sc_hd__clkbuf_1
X_544_ clknet_3_4__leaf_clk _062_ VGND VGND VPWR VPWR registers\[7\]\[6\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_28_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_260_ registers\[2\]\[3\] registers\[3\]\[3\] _072_ VGND VGND VPWR VPWR _088_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_389_ _182_ VGND VGND VPWR VPWR _021_ sky130_fd_sc_hd__clkbuf_1
X_458_ net57 net13 _214_ VGND VGND VPWR VPWR _220_ sky130_fd_sc_hd__mux2_1
X_527_ clknet_3_5__leaf_clk _045_ VGND VGND VPWR VPWR registers\[0\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_243_ _069_ _071_ _073_ _067_ net6 VGND VGND VPWR VPWR _074_ sky130_fd_sc_hd__a221o_1
X_312_ registers\[1\]\[3\] _116_ VGND VGND VPWR VPWR _132_ sky130_fd_sc_hd__or2b_1
Xinput18 writeReg[2] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_TAPCELL_ROW_30_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold7 registers\[2\]\[0\] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_491_ clknet_3_0__leaf_clk _009_ VGND VGND VPWR VPWR registers\[5\]\[1\] sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_543_ clknet_3_6__leaf_clk _061_ VGND VGND VPWR VPWR registers\[7\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_474_ net81 net12 _224_ VGND VGND VPWR VPWR _229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_526_ clknet_3_7__leaf_clk _044_ VGND VGND VPWR VPWR registers\[0\]\[4\] sky130_fd_sc_hd__dfxtp_1
X_388_ net80 net13 _176_ VGND VGND VPWR VPWR _182_ sky130_fd_sc_hd__mux2_1
X_457_ _219_ VGND VGND VPWR VPWR _052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_311_ registers\[4\]\[3\] registers\[5\]\[3\] registers\[6\]\[3\] registers\[7\]\[3\]
+ _111_ _112_ VGND VGND VPWR VPWR _131_ sky130_fd_sc_hd__mux4_1
X_242_ registers\[2\]\[0\] registers\[3\]\[0\] _072_ VGND VGND VPWR VPWR _073_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_30_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_509_ clknet_3_3__leaf_clk _027_ VGND VGND VPWR VPWR registers\[3\]\[3\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_2_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_5_Left_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold8 registers\[6\]\[5\] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_7 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_490_ clknet_3_2__leaf_clk _008_ VGND VGND VPWR VPWR registers\[5\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_473_ _228_ VGND VGND VPWR VPWR _059_ sky130_fd_sc_hd__clkbuf_1
X_542_ clknet_3_6__leaf_clk _060_ VGND VGND VPWR VPWR registers\[7\]\[4\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_387_ _181_ VGND VGND VPWR VPWR _020_ sky130_fd_sc_hd__clkbuf_1
X_456_ net63 net12 _214_ VGND VGND VPWR VPWR _219_ sky130_fd_sc_hd__mux2_1
X_525_ clknet_3_6__leaf_clk _043_ VGND VGND VPWR VPWR registers\[0\]\[3\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_310_ _110_ _126_ _130_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__o21a_1
X_439_ net12 net93 _205_ VGND VGND VPWR VPWR _210_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_15_110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_241_ net4 VGND VGND VPWR VPWR _072_ sky130_fd_sc_hd__clkbuf_4
X_508_ clknet_3_0__leaf_clk _026_ VGND VGND VPWR VPWR registers\[3\]\[2\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_30_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_21_Left_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_12_102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold9 registers\[2\]\[1\] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_15_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_541_ clknet_3_3__leaf_clk _059_ VGND VGND VPWR VPWR registers\[7\]\[3\] sky130_fd_sc_hd__dfxtp_1
X_472_ net78 net11 _224_ VGND VGND VPWR VPWR _228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_386_ net39 net12 _176_ VGND VGND VPWR VPWR _181_ sky130_fd_sc_hd__mux2_1
X_455_ _218_ VGND VGND VPWR VPWR _051_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_2_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_524_ clknet_3_1__leaf_clk _042_ VGND VGND VPWR VPWR registers\[0\]\[2\] sky130_fd_sc_hd__dfxtp_1
X_240_ registers\[0\]\[0\] _070_ _066_ VGND VGND VPWR VPWR _071_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_30_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_369_ net71 net12 _167_ VGND VGND VPWR VPWR _172_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_438_ _209_ VGND VGND VPWR VPWR _043_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_15_111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_507_ clknet_3_2__leaf_clk _025_ VGND VGND VPWR VPWR registers\[3\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_12_103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_471_ _227_ VGND VGND VPWR VPWR _058_ sky130_fd_sc_hd__clkbuf_1
X_540_ clknet_3_0__leaf_clk _058_ VGND VGND VPWR VPWR registers\[7\]\[2\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_385_ _180_ VGND VGND VPWR VPWR _019_ sky130_fd_sc_hd__clkbuf_1
X_454_ net58 net11 _214_ VGND VGND VPWR VPWR _218_ sky130_fd_sc_hd__mux2_1
X_523_ clknet_3_3__leaf_clk _041_ VGND VGND VPWR VPWR registers\[0\]\[1\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_2_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_368_ _171_ VGND VGND VPWR VPWR _011_ sky130_fd_sc_hd__clkbuf_1
X_506_ clknet_3_2__leaf_clk _024_ VGND VGND VPWR VPWR registers\[3\]\[0\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_15_112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_437_ net11 net97 _205_ VGND VGND VPWR VPWR _209_ sky130_fd_sc_hd__mux2_1
X_299_ registers\[4\]\[1\] registers\[5\]\[1\] registers\[6\]\[1\] registers\[7\]\[1\]
+ _111_ _113_ VGND VGND VPWR VPWR _121_ sky130_fd_sc_hd__mux4_1
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_470_ net59 net10 _224_ VGND VGND VPWR VPWR _227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_384_ net68 net11 _176_ VGND VGND VPWR VPWR _180_ sky130_fd_sc_hd__mux2_1
X_522_ clknet_3_3__leaf_clk _040_ VGND VGND VPWR VPWR registers\[0\]\[0\] sky130_fd_sc_hd__dfxtp_1
XFILLER_0_8_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_453_ _217_ VGND VGND VPWR VPWR _050_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_18_121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_367_ net62 net11 _167_ VGND VGND VPWR VPWR _171_ sky130_fd_sc_hd__mux2_1
X_298_ _110_ _114_ _120_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__o21a_1
X_505_ clknet_3_4__leaf_clk _023_ VGND VGND VPWR VPWR registers\[4\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_436_ _208_ VGND VGND VPWR VPWR _042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_25_Left_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_419_ net77 net11 _195_ VGND VGND VPWR VPWR _199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_1 readReg2[1] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_383_ _179_ VGND VGND VPWR VPWR _018_ sky130_fd_sc_hd__clkbuf_1
X_521_ clknet_3_5__leaf_clk _039_ VGND VGND VPWR VPWR registers\[2\]\[7\] sky130_fd_sc_hd__dfxtp_1
X_452_ net89 net10 _214_ VGND VGND VPWR VPWR _217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_297_ _115_ _117_ _119_ _113_ net3 VGND VGND VPWR VPWR _120_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_504_ clknet_3_5__leaf_clk _022_ VGND VGND VPWR VPWR registers\[4\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_366_ _170_ VGND VGND VPWR VPWR _010_ sky130_fd_sc_hd__clkbuf_1
X_435_ net10 net95 _205_ VGND VGND VPWR VPWR _208_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_0_Left_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_349_ net37 net11 _157_ VGND VGND VPWR VPWR _161_ sky130_fd_sc_hd__mux2_1
X_418_ _198_ VGND VGND VPWR VPWR _034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold60 registers\[0\]\[1\] VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlygate4sd3_1
X_520_ clknet_3_5__leaf_clk _038_ VGND VGND VPWR VPWR registers\[2\]\[6\] sky130_fd_sc_hd__dfxtp_1
X_451_ _216_ VGND VGND VPWR VPWR _049_ sky130_fd_sc_hd__clkbuf_1
X_382_ net67 net10 _176_ VGND VGND VPWR VPWR _179_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_24_137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_503_ clknet_3_7__leaf_clk _021_ VGND VGND VPWR VPWR registers\[4\]\[5\] sky130_fd_sc_hd__dfxtp_1
X_296_ registers\[2\]\[0\] registers\[3\]\[0\] _118_ VGND VGND VPWR VPWR _119_ sky130_fd_sc_hd__mux2_1
X_434_ _207_ VGND VGND VPWR VPWR _041_ sky130_fd_sc_hd__clkbuf_1
X_365_ net46 net10 _167_ VGND VGND VPWR VPWR _170_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_21_129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_348_ _160_ VGND VGND VPWR VPWR _002_ sky130_fd_sc_hd__clkbuf_1
X_417_ net47 net10 _195_ VGND VGND VPWR VPWR _198_ sky130_fd_sc_hd__mux2_1
X_279_ _101_ _102_ _103_ _067_ net6 VGND VGND VPWR VPWR _104_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold50 registers\[4\]\[0\] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold61 registers\[0\]\[2\] VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_TAPCELL_ROW_27_146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_450_ net40 net9 _214_ VGND VGND VPWR VPWR _216_ sky130_fd_sc_hd__mux2_1
X_381_ _178_ VGND VGND VPWR VPWR _017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_502_ clknet_3_7__leaf_clk _020_ VGND VGND VPWR VPWR registers\[4\]\[4\] sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_24_138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_433_ net9 net94 _205_ VGND VGND VPWR VPWR _207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_295_ net1 VGND VGND VPWR VPWR _118_ sky130_fd_sc_hd__clkbuf_4
X_364_ _169_ VGND VGND VPWR VPWR _009_ sky130_fd_sc_hd__clkbuf_1
X_416_ _197_ VGND VGND VPWR VPWR _033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_347_ net65 net10 _157_ VGND VGND VPWR VPWR _160_ sky130_fd_sc_hd__mux2_1
X_278_ registers\[2\]\[6\] registers\[3\]\[6\] net4 VGND VGND VPWR VPWR _103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xhold51 registers\[3\]\[3\] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 registers\[0\]\[6\] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlygate4sd3_1
Xhold40 registers\[5\]\[6\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_21_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_16_Left_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput30 net30 VGND VGND VPWR VPWR readData2[3] sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_27_147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_380_ net64 net9 _176_ VGND VGND VPWR VPWR _178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
.ends

