magic
tech sky130A
magscale 1 2
timestamp 1748200543
<< nwell >>
rect 1066 2159 18162 19078
<< obsli1 >>
rect 1104 2159 18124 19057
<< obsm1 >>
rect 842 2128 18124 19088
<< metal2 >>
rect 9034 20613 9090 21413
rect 9678 20613 9734 21413
rect 10322 20613 10378 21413
rect 12898 20613 12954 21413
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
<< obsm2 >>
rect 846 20557 8978 20754
rect 9146 20557 9622 20754
rect 9790 20557 10266 20754
rect 10434 20557 12842 20754
rect 13010 20557 17830 20754
rect 846 856 17830 20557
rect 846 800 3826 856
rect 3994 800 6402 856
rect 6570 800 7046 856
rect 7214 800 8334 856
rect 8502 800 8978 856
rect 9146 800 9622 856
rect 9790 800 10266 856
rect 10434 800 10910 856
rect 11078 800 11554 856
rect 11722 800 12198 856
rect 12366 800 17830 856
<< metal3 >>
rect 0 17688 800 17808
rect 0 16328 800 16448
rect 18469 15648 19269 15768
rect 0 14968 800 15088
rect 18469 14968 19269 15088
rect 0 14288 800 14408
rect 18469 14288 19269 14408
rect 0 12928 800 13048
rect 18469 12928 19269 13048
rect 0 12248 800 12368
rect 0 10888 800 11008
rect 0 10208 800 10328
rect 18469 10208 19269 10328
rect 0 9528 800 9648
rect 18469 8168 19269 8288
rect 18469 7488 19269 7608
rect 18469 6808 19269 6928
rect 18469 6128 19269 6248
rect 18469 5448 19269 5568
rect 18469 4768 19269 4888
rect 18469 3408 19269 3528
<< obsm3 >>
rect 798 17888 18469 19073
rect 880 17608 18469 17888
rect 798 16528 18469 17608
rect 880 16248 18469 16528
rect 798 15848 18469 16248
rect 798 15568 18389 15848
rect 798 15168 18469 15568
rect 880 14888 18389 15168
rect 798 14488 18469 14888
rect 880 14208 18389 14488
rect 798 13128 18469 14208
rect 880 12848 18389 13128
rect 798 12448 18469 12848
rect 880 12168 18469 12448
rect 798 11088 18469 12168
rect 880 10808 18469 11088
rect 798 10408 18469 10808
rect 880 10128 18389 10408
rect 798 9728 18469 10128
rect 880 9448 18469 9728
rect 798 8368 18469 9448
rect 798 8088 18389 8368
rect 798 7688 18469 8088
rect 798 7408 18389 7688
rect 798 7008 18469 7408
rect 798 6728 18389 7008
rect 798 6328 18469 6728
rect 798 6048 18389 6328
rect 798 5648 18469 6048
rect 798 5368 18389 5648
rect 798 4968 18469 5368
rect 798 4688 18389 4968
rect 798 3608 18469 4688
rect 798 3328 18389 3608
rect 798 2143 18469 3328
<< metal4 >>
rect 3071 2128 3391 19088
rect 3731 2128 4051 19088
rect 7326 2128 7646 19088
rect 7986 2128 8306 19088
rect 11581 2128 11901 19088
rect 12241 2128 12561 19088
rect 15836 2128 16156 19088
rect 16496 2128 16816 19088
<< obsm4 >>
rect 3555 5747 3651 17781
rect 4131 5747 7246 17781
rect 7726 5747 7906 17781
rect 8386 5747 11501 17781
rect 11981 5747 12161 17781
rect 12641 5747 14477 17781
<< metal5 >>
rect 1056 17432 18172 17752
rect 1056 16772 18172 17092
rect 1056 13216 18172 13536
rect 1056 12556 18172 12876
rect 1056 9000 18172 9320
rect 1056 8340 18172 8660
rect 1056 4784 18172 5104
rect 1056 4124 18172 4444
<< labels >>
rlabel metal4 s 3731 2128 4051 19088 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 7986 2128 8306 19088 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12241 2128 12561 19088 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 16496 2128 16816 19088 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 4784 18172 5104 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 9000 18172 9320 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 13216 18172 13536 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 17432 18172 17752 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 3071 2128 3391 19088 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 7326 2128 7646 19088 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11581 2128 11901 19088 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 15836 2128 16156 19088 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 4124 18172 4444 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 8340 18172 8660 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 12556 18172 12876 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 16772 18172 17092 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 17688 800 17808 6 clk
port 3 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 readData1[0]
port 4 nsew signal output
rlabel metal3 s 0 9528 800 9648 6 readData1[1]
port 5 nsew signal output
rlabel metal2 s 6458 0 6514 800 6 readData1[2]
port 6 nsew signal output
rlabel metal2 s 9678 20613 9734 21413 6 readData1[3]
port 7 nsew signal output
rlabel metal3 s 18469 15648 19269 15768 6 readData1[4]
port 8 nsew signal output
rlabel metal2 s 12898 20613 12954 21413 6 readData1[5]
port 9 nsew signal output
rlabel metal3 s 18469 5448 19269 5568 6 readData1[6]
port 10 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 readData1[7]
port 11 nsew signal output
rlabel metal3 s 0 14288 800 14408 6 readData2[0]
port 12 nsew signal output
rlabel metal3 s 0 10208 800 10328 6 readData2[1]
port 13 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 readData2[2]
port 14 nsew signal output
rlabel metal2 s 10322 20613 10378 21413 6 readData2[3]
port 15 nsew signal output
rlabel metal3 s 18469 14968 19269 15088 6 readData2[4]
port 16 nsew signal output
rlabel metal3 s 18469 14288 19269 14408 6 readData2[5]
port 17 nsew signal output
rlabel metal3 s 18469 4768 19269 4888 6 readData2[6]
port 18 nsew signal output
rlabel metal2 s 10966 0 11022 800 6 readData2[7]
port 19 nsew signal output
rlabel metal3 s 18469 6128 19269 6248 6 readReg1[0]
port 20 nsew signal input
rlabel metal3 s 18469 7488 19269 7608 6 readReg1[1]
port 21 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 readReg1[2]
port 22 nsew signal input
rlabel metal3 s 18469 6808 19269 6928 6 readReg2[0]
port 23 nsew signal input
rlabel metal3 s 18469 8168 19269 8288 6 readReg2[1]
port 24 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 readReg2[2]
port 25 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 regWrite
port 26 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 writeData[0]
port 27 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 writeData[1]
port 28 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 writeData[2]
port 29 nsew signal input
rlabel metal2 s 9034 20613 9090 21413 6 writeData[3]
port 30 nsew signal input
rlabel metal3 s 18469 12928 19269 13048 6 writeData[4]
port 31 nsew signal input
rlabel metal3 s 18469 10208 19269 10328 6 writeData[5]
port 32 nsew signal input
rlabel metal3 s 18469 3408 19269 3528 6 writeData[6]
port 33 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 writeData[7]
port 34 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 writeReg[0]
port 35 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 writeReg[1]
port 36 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 writeReg[2]
port 37 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 19269 21413
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1201656
string GDS_FILE /openlane/designs/register_file/runs/RUN_2025.05.25_19.14.43/results/signoff/register_file.magic.gds
string GDS_START 190606
<< end >>

