VERSION 5.8 ;
SITE CoreSite ;
MACRO INVX1 ;
