magic
tech sky130A
magscale 1 2
timestamp 1748200542
<< viali >>
rect 10057 18921 10091 18955
rect 12633 18921 12667 18955
rect 7113 18717 7147 18751
rect 7481 18717 7515 18751
rect 8401 18717 8435 18751
rect 8677 18717 8711 18751
rect 9505 18717 9539 18751
rect 10793 18717 10827 18751
rect 11161 18717 11195 18751
rect 12173 18717 12207 18751
rect 13461 18717 13495 18751
rect 13829 18717 13863 18751
rect 8493 18649 8527 18683
rect 9781 18649 9815 18683
rect 12725 18649 12759 18683
rect 6929 18581 6963 18615
rect 7665 18581 7699 18615
rect 7757 18581 7791 18615
rect 8953 18581 8987 18615
rect 10241 18581 10275 18615
rect 11345 18581 11379 18615
rect 11529 18581 11563 18615
rect 12909 18581 12943 18615
rect 13645 18581 13679 18615
rect 9321 18377 9355 18411
rect 9505 18377 9539 18411
rect 13093 18377 13127 18411
rect 8186 18309 8220 18343
rect 9781 18309 9815 18343
rect 13544 18309 13578 18343
rect 6469 18241 6503 18275
rect 6736 18241 6770 18275
rect 9965 18241 9999 18275
rect 10232 18241 10266 18275
rect 11713 18241 11747 18275
rect 11969 18241 12003 18275
rect 13277 18241 13311 18275
rect 15669 18241 15703 18275
rect 7941 18173 7975 18207
rect 15301 18173 15335 18207
rect 14657 18105 14691 18139
rect 7849 18037 7883 18071
rect 11345 18037 11379 18071
rect 14749 18037 14783 18071
rect 15485 18037 15519 18071
rect 7205 17833 7239 17867
rect 8033 17833 8067 17867
rect 10517 17833 10551 17867
rect 10701 17833 10735 17867
rect 12173 17833 12207 17867
rect 13921 17833 13955 17867
rect 14289 17833 14323 17867
rect 6745 17697 6779 17731
rect 6929 17697 6963 17731
rect 7849 17697 7883 17731
rect 8677 17697 8711 17731
rect 11529 17697 11563 17731
rect 12725 17697 12759 17731
rect 13277 17697 13311 17731
rect 16313 17697 16347 17731
rect 4721 17629 4755 17663
rect 5089 17629 5123 17663
rect 5641 17629 5675 17663
rect 7573 17629 7607 17663
rect 9137 17629 9171 17663
rect 10885 17629 10919 17663
rect 11345 17629 11379 17663
rect 12541 17629 12575 17663
rect 15402 17629 15436 17663
rect 15669 17629 15703 17663
rect 6193 17561 6227 17595
rect 6653 17561 6687 17595
rect 8401 17561 8435 17595
rect 9404 17561 9438 17595
rect 13553 17561 13587 17595
rect 4169 17493 4203 17527
rect 4905 17493 4939 17527
rect 6285 17493 6319 17527
rect 7665 17493 7699 17527
rect 8493 17493 8527 17527
rect 10977 17493 11011 17527
rect 11437 17493 11471 17527
rect 12633 17493 12667 17527
rect 13461 17493 13495 17527
rect 15761 17493 15795 17527
rect 3985 17289 4019 17323
rect 6193 17289 6227 17323
rect 9781 17289 9815 17323
rect 10241 17289 10275 17323
rect 14473 17289 14507 17323
rect 14565 17289 14599 17323
rect 14933 17289 14967 17323
rect 4528 17221 4562 17255
rect 2872 17153 2906 17187
rect 6009 17153 6043 17187
rect 7490 17153 7524 17187
rect 9689 17153 9723 17187
rect 10425 17153 10459 17187
rect 2605 17085 2639 17119
rect 4261 17085 4295 17119
rect 7757 17085 7791 17119
rect 9505 17085 9539 17119
rect 11345 17085 11379 17119
rect 14289 17085 14323 17119
rect 6377 17017 6411 17051
rect 10149 17017 10183 17051
rect 5641 16949 5675 16983
rect 10701 16949 10735 16983
rect 2973 16745 3007 16779
rect 4721 16745 4755 16779
rect 11713 16745 11747 16779
rect 8309 16677 8343 16711
rect 15485 16677 15519 16711
rect 1685 16609 1719 16643
rect 4445 16609 4479 16643
rect 5181 16609 5215 16643
rect 5365 16609 5399 16643
rect 6101 16609 6135 16643
rect 9505 16609 9539 16643
rect 10333 16609 10367 16643
rect 11897 16609 11931 16643
rect 12541 16609 12575 16643
rect 12934 16609 12968 16643
rect 13093 16609 13127 16643
rect 13737 16609 13771 16643
rect 15577 16609 15611 16643
rect 3157 16541 3191 16575
rect 4169 16541 4203 16575
rect 4261 16541 4295 16575
rect 6929 16541 6963 16575
rect 12081 16541 12115 16575
rect 12817 16541 12851 16575
rect 15301 16541 15335 16575
rect 17601 16541 17635 16575
rect 1501 16473 1535 16507
rect 5089 16473 5123 16507
rect 5549 16473 5583 16507
rect 7196 16473 7230 16507
rect 10600 16473 10634 16507
rect 15822 16473 15856 16507
rect 3801 16405 3835 16439
rect 8953 16405 8987 16439
rect 16957 16405 16991 16439
rect 17049 16405 17083 16439
rect 7205 16201 7239 16235
rect 7849 16201 7883 16235
rect 10977 16201 11011 16235
rect 11345 16201 11379 16235
rect 11529 16201 11563 16235
rect 15485 16201 15519 16235
rect 15853 16201 15887 16235
rect 10885 16133 10919 16167
rect 15945 16133 15979 16167
rect 3157 16065 3191 16099
rect 3424 16065 3458 16099
rect 5181 16065 5215 16099
rect 7389 16065 7423 16099
rect 8585 16065 8619 16099
rect 9622 16065 9656 16099
rect 11713 16065 11747 16099
rect 11897 16065 11931 16099
rect 12081 16065 12115 16099
rect 12817 16065 12851 16099
rect 12934 16065 12968 16099
rect 17509 16065 17543 16099
rect 7941 15997 7975 16031
rect 8033 15997 8067 16031
rect 8769 15997 8803 16031
rect 9505 15997 9539 16031
rect 9781 15997 9815 16031
rect 10793 15997 10827 16031
rect 13093 15997 13127 16031
rect 16037 15997 16071 16031
rect 17233 15997 17267 16031
rect 4537 15929 4571 15963
rect 7481 15929 7515 15963
rect 9229 15929 9263 15963
rect 12541 15929 12575 15963
rect 4629 15861 4663 15895
rect 10425 15861 10459 15895
rect 13737 15861 13771 15895
rect 16681 15861 16715 15895
rect 17693 15861 17727 15895
rect 3433 15657 3467 15691
rect 3801 15589 3835 15623
rect 4261 15521 4295 15555
rect 4445 15521 4479 15555
rect 5457 15521 5491 15555
rect 5850 15521 5884 15555
rect 6009 15521 6043 15555
rect 8953 15521 8987 15555
rect 9137 15521 9171 15555
rect 9597 15521 9631 15555
rect 9990 15521 10024 15555
rect 10149 15521 10183 15555
rect 15301 15521 15335 15555
rect 16037 15521 16071 15555
rect 1685 15453 1719 15487
rect 3617 15453 3651 15487
rect 4169 15453 4203 15487
rect 4813 15453 4847 15487
rect 4997 15453 5031 15487
rect 5733 15453 5767 15487
rect 7481 15453 7515 15487
rect 9873 15453 9907 15487
rect 13185 15453 13219 15487
rect 14749 15453 14783 15487
rect 14887 15453 14921 15487
rect 15025 15453 15059 15487
rect 15761 15453 15795 15487
rect 15945 15453 15979 15487
rect 17509 15453 17543 15487
rect 16304 15385 16338 15419
rect 1501 15317 1535 15351
rect 6653 15317 6687 15351
rect 7297 15317 7331 15351
rect 10793 15317 10827 15351
rect 12541 15317 12575 15351
rect 14105 15317 14139 15351
rect 17417 15317 17451 15351
rect 17693 15317 17727 15351
rect 9965 15113 9999 15147
rect 10517 15113 10551 15147
rect 11345 15113 11379 15147
rect 12909 15113 12943 15147
rect 15853 15113 15887 15147
rect 16221 15113 16255 15147
rect 16313 15113 16347 15147
rect 7196 15045 7230 15079
rect 11774 15045 11808 15079
rect 1768 14977 1802 15011
rect 4353 14977 4387 15011
rect 5273 14977 5307 15011
rect 5390 14977 5424 15011
rect 6561 14977 6595 15011
rect 6745 14977 6779 15011
rect 6837 14977 6871 15011
rect 9321 14977 9355 15011
rect 10149 14977 10183 15011
rect 10333 14977 10367 15011
rect 10701 14977 10735 15011
rect 10885 14977 10919 15011
rect 10977 14977 11011 15011
rect 11161 14977 11195 15011
rect 13896 14977 13930 15011
rect 16497 14977 16531 15011
rect 17785 14977 17819 15011
rect 1501 14909 1535 14943
rect 3525 14909 3559 14943
rect 4537 14909 4571 14943
rect 5549 14909 5583 14943
rect 6929 14909 6963 14943
rect 8953 14909 8987 14943
rect 10425 14909 10459 14943
rect 11529 14909 11563 14943
rect 13737 14909 13771 14943
rect 14013 14909 14047 14943
rect 14749 14909 14783 14943
rect 14933 14909 14967 14943
rect 15669 14909 15703 14943
rect 15761 14909 15795 14943
rect 17417 14909 17451 14943
rect 2973 14841 3007 14875
rect 4997 14841 5031 14875
rect 8309 14841 8343 14875
rect 14289 14841 14323 14875
rect 2881 14773 2915 14807
rect 6193 14773 6227 14807
rect 6377 14773 6411 14807
rect 8401 14773 8435 14807
rect 9137 14773 9171 14807
rect 13093 14773 13127 14807
rect 16865 14773 16899 14807
rect 17601 14773 17635 14807
rect 1961 14569 1995 14603
rect 6101 14569 6135 14603
rect 6469 14569 6503 14603
rect 10333 14569 10367 14603
rect 14105 14569 14139 14603
rect 14473 14569 14507 14603
rect 14749 14569 14783 14603
rect 15117 14569 15151 14603
rect 16313 14569 16347 14603
rect 1501 14501 1535 14535
rect 16405 14501 16439 14535
rect 2881 14433 2915 14467
rect 6561 14433 6595 14467
rect 10977 14433 11011 14467
rect 11897 14433 11931 14467
rect 14565 14433 14599 14467
rect 14657 14433 14691 14467
rect 15761 14433 15795 14467
rect 1685 14365 1719 14399
rect 2145 14365 2179 14399
rect 2697 14365 2731 14399
rect 6285 14365 6319 14399
rect 8953 14365 8987 14399
rect 9220 14365 9254 14399
rect 11621 14365 11655 14399
rect 14289 14365 14323 14399
rect 14933 14365 14967 14399
rect 17518 14365 17552 14399
rect 17785 14365 17819 14399
rect 7021 14297 7055 14331
rect 8769 14297 8803 14331
rect 13645 14297 13679 14331
rect 15853 14297 15887 14331
rect 15945 14297 15979 14331
rect 2329 14229 2363 14263
rect 2789 14229 2823 14263
rect 10425 14229 10459 14263
rect 6377 14025 6411 14059
rect 7481 14025 7515 14059
rect 7849 14025 7883 14059
rect 9321 14025 9355 14059
rect 10057 14025 10091 14059
rect 10149 14025 10183 14059
rect 11621 14025 11655 14059
rect 11989 14025 12023 14059
rect 14749 14025 14783 14059
rect 15117 14025 15151 14059
rect 15945 14025 15979 14059
rect 16957 14025 16991 14059
rect 4353 13957 4387 13991
rect 6745 13957 6779 13991
rect 8953 13957 8987 13991
rect 12081 13957 12115 13991
rect 16037 13957 16071 13991
rect 1961 13889 1995 13923
rect 5273 13889 5307 13923
rect 6515 13889 6549 13923
rect 6653 13889 6687 13923
rect 6928 13889 6962 13923
rect 7021 13889 7055 13923
rect 7941 13889 7975 13923
rect 12633 13889 12667 13923
rect 13185 13889 13219 13923
rect 13277 13889 13311 13923
rect 13461 13889 13495 13923
rect 14197 13889 14231 13923
rect 14289 13889 14323 13923
rect 14473 13889 14507 13923
rect 16773 13889 16807 13923
rect 17693 13889 17727 13923
rect 3341 13821 3375 13855
rect 5733 13821 5767 13855
rect 8033 13821 8067 13855
rect 8677 13821 8711 13855
rect 8861 13821 8895 13855
rect 10333 13821 10367 13855
rect 12173 13821 12207 13855
rect 15209 13821 15243 13855
rect 15301 13821 15335 13855
rect 16129 13821 16163 13855
rect 13645 13753 13679 13787
rect 1777 13685 1811 13719
rect 2697 13685 2731 13719
rect 5549 13685 5583 13719
rect 9689 13685 9723 13719
rect 12449 13685 12483 13719
rect 14657 13685 14691 13719
rect 15577 13685 15611 13719
rect 17141 13685 17175 13719
rect 10425 13481 10459 13515
rect 16037 13481 16071 13515
rect 2789 13413 2823 13447
rect 10333 13413 10367 13447
rect 12725 13413 12759 13447
rect 3065 13345 3099 13379
rect 3157 13345 3191 13379
rect 4261 13345 4295 13379
rect 9781 13345 9815 13379
rect 11345 13345 11379 13379
rect 13369 13345 13403 13379
rect 16773 13345 16807 13379
rect 1409 13277 1443 13311
rect 1676 13277 1710 13311
rect 3249 13277 3283 13311
rect 6009 13277 6043 13311
rect 6561 13277 6595 13311
rect 6837 13277 6871 13311
rect 7021 13277 7055 13311
rect 9873 13277 9907 13311
rect 10604 13277 10638 13311
rect 10701 13277 10735 13311
rect 10793 13277 10827 13311
rect 10976 13277 11010 13311
rect 11069 13277 11103 13311
rect 11612 13277 11646 13311
rect 14749 13277 14783 13311
rect 16865 13277 16899 13311
rect 16957 13277 16991 13311
rect 17509 13277 17543 13311
rect 9965 13209 9999 13243
rect 14473 13209 14507 13243
rect 17693 13209 17727 13243
rect 3617 13141 3651 13175
rect 6377 13141 6411 13175
rect 12817 13141 12851 13175
rect 17325 13141 17359 13175
rect 2145 12937 2179 12971
rect 2513 12937 2547 12971
rect 3249 12937 3283 12971
rect 5181 12937 5215 12971
rect 6193 12937 6227 12971
rect 6837 12937 6871 12971
rect 10425 12937 10459 12971
rect 12173 12937 12207 12971
rect 12633 12937 12667 12971
rect 13921 12937 13955 12971
rect 14657 12937 14691 12971
rect 17417 12937 17451 12971
rect 1501 12869 1535 12903
rect 3341 12869 3375 12903
rect 5825 12869 5859 12903
rect 7174 12869 7208 12903
rect 10057 12869 10091 12903
rect 12265 12869 12299 12903
rect 13553 12869 13587 12903
rect 14289 12869 14323 12903
rect 16252 12869 16286 12903
rect 3801 12801 3835 12835
rect 4068 12801 4102 12835
rect 5549 12801 5583 12835
rect 5697 12801 5731 12835
rect 5917 12801 5951 12835
rect 6055 12801 6089 12835
rect 6653 12801 6687 12835
rect 9229 12801 9263 12835
rect 9781 12801 9815 12835
rect 9929 12801 9963 12835
rect 10149 12801 10183 12835
rect 10287 12801 10321 12835
rect 10701 12801 10735 12835
rect 10885 12801 10919 12835
rect 11161 12801 11195 12835
rect 11345 12801 11379 12835
rect 12725 12801 12759 12835
rect 13277 12801 13311 12835
rect 13370 12801 13404 12835
rect 13645 12801 13679 12835
rect 13742 12801 13776 12835
rect 14013 12801 14047 12835
rect 14161 12801 14195 12835
rect 14381 12801 14415 12835
rect 14478 12801 14512 12835
rect 17601 12801 17635 12835
rect 2605 12733 2639 12767
rect 2697 12733 2731 12767
rect 3065 12733 3099 12767
rect 6929 12733 6963 12767
rect 8953 12733 8987 12767
rect 9689 12733 9723 12767
rect 12081 12733 12115 12767
rect 13185 12733 13219 12767
rect 16497 12733 16531 12767
rect 17233 12733 17267 12767
rect 1777 12597 1811 12631
rect 3709 12597 3743 12631
rect 8309 12597 8343 12631
rect 8401 12597 8435 12631
rect 9413 12597 9447 12631
rect 13001 12597 13035 12631
rect 15117 12597 15151 12631
rect 16681 12597 16715 12631
rect 3985 12393 4019 12427
rect 5825 12393 5859 12427
rect 6009 12393 6043 12427
rect 6377 12393 6411 12427
rect 7113 12393 7147 12427
rect 9505 12393 9539 12427
rect 10701 12393 10735 12427
rect 13001 12393 13035 12427
rect 14289 12393 14323 12427
rect 16313 12393 16347 12427
rect 16405 12393 16439 12427
rect 13277 12325 13311 12359
rect 4813 12257 4847 12291
rect 5733 12257 5767 12291
rect 7573 12257 7607 12291
rect 7757 12257 7791 12291
rect 9873 12257 9907 12291
rect 15669 12257 15703 12291
rect 15853 12257 15887 12291
rect 1501 12189 1535 12223
rect 2145 12189 2179 12223
rect 3341 12189 3375 12223
rect 4169 12189 4203 12223
rect 6285 12189 6319 12223
rect 6561 12189 6595 12223
rect 6837 12189 6871 12223
rect 7021 12189 7055 12223
rect 8401 12189 8435 12223
rect 8953 12189 8987 12223
rect 9413 12189 9447 12223
rect 10885 12189 10919 12223
rect 11161 12189 11195 12223
rect 11345 12189 11379 12223
rect 12817 12189 12851 12223
rect 14473 12189 14507 12223
rect 14749 12189 14783 12223
rect 14933 12189 14967 12223
rect 17785 12189 17819 12223
rect 4629 12121 4663 12155
rect 5089 12121 5123 12155
rect 15945 12121 15979 12155
rect 17540 12121 17574 12155
rect 1777 12053 1811 12087
rect 1961 12053 1995 12087
rect 2789 12053 2823 12087
rect 4261 12053 4295 12087
rect 4721 12053 4755 12087
rect 7481 12053 7515 12087
rect 8493 12053 8527 12087
rect 9045 12053 9079 12087
rect 8769 11849 8803 11883
rect 14105 11849 14139 11883
rect 17693 11849 17727 11883
rect 9229 11781 9263 11815
rect 1860 11713 1894 11747
rect 3617 11713 3651 11747
rect 3884 11713 3918 11747
rect 6561 11713 6595 11747
rect 6837 11713 6871 11747
rect 7021 11713 7055 11747
rect 8677 11713 8711 11747
rect 9137 11713 9171 11747
rect 9597 11713 9631 11747
rect 11713 11713 11747 11747
rect 12633 11713 12667 11747
rect 13553 11713 13587 11747
rect 13829 11713 13863 11747
rect 14013 11713 14047 11747
rect 14289 11713 14323 11747
rect 14565 11713 14599 11747
rect 14749 11713 14783 11747
rect 15577 11713 15611 11747
rect 16497 11713 16531 11747
rect 17049 11713 17083 11747
rect 17509 11713 17543 11747
rect 1593 11645 1627 11679
rect 5641 11645 5675 11679
rect 9321 11645 9355 11679
rect 10149 11645 10183 11679
rect 15945 11645 15979 11679
rect 17141 11645 17175 11679
rect 17233 11645 17267 11679
rect 5089 11577 5123 11611
rect 13093 11577 13127 11611
rect 16681 11577 16715 11611
rect 2973 11509 3007 11543
rect 4997 11509 5031 11543
rect 6377 11509 6411 11543
rect 8493 11509 8527 11543
rect 11529 11509 11563 11543
rect 12725 11509 12759 11543
rect 13369 11509 13403 11543
rect 15761 11509 15795 11543
rect 2053 11305 2087 11339
rect 3985 11305 4019 11339
rect 5365 11305 5399 11339
rect 4261 11237 4295 11271
rect 16405 11237 16439 11271
rect 2605 11169 2639 11203
rect 2973 11169 3007 11203
rect 4813 11169 4847 11203
rect 7849 11169 7883 11203
rect 15301 11169 15335 11203
rect 16129 11169 16163 11203
rect 1961 11101 1995 11135
rect 2421 11101 2455 11135
rect 4169 11101 4203 11135
rect 4629 11101 4663 11135
rect 4721 11101 4755 11135
rect 5089 11101 5123 11135
rect 5641 11101 5675 11135
rect 5789 11101 5823 11135
rect 6147 11101 6181 11135
rect 6469 11101 6503 11135
rect 6653 11101 6687 11135
rect 6929 11101 6963 11135
rect 7113 11101 7147 11135
rect 8677 11101 8711 11135
rect 9505 11101 9539 11135
rect 9781 11101 9815 11135
rect 11253 11101 11287 11135
rect 11520 11101 11554 11135
rect 13277 11101 13311 11135
rect 15117 11101 15151 11135
rect 15945 11101 15979 11135
rect 17785 11101 17819 11135
rect 1501 11033 1535 11067
rect 1685 11033 1719 11067
rect 5917 11033 5951 11067
rect 6009 11033 6043 11067
rect 7665 11033 7699 11067
rect 7757 11033 7791 11067
rect 8125 11033 8159 11067
rect 10026 11033 10060 11067
rect 12725 11033 12759 11067
rect 15209 11033 15243 11067
rect 17518 11033 17552 11067
rect 1777 10965 1811 10999
rect 2513 10965 2547 10999
rect 3157 10965 3191 10999
rect 3249 10965 3283 10999
rect 3617 10965 3651 10999
rect 5549 10965 5583 10999
rect 6285 10965 6319 10999
rect 7297 10965 7331 10999
rect 9689 10965 9723 10999
rect 11161 10965 11195 10999
rect 12633 10965 12667 10999
rect 14749 10965 14783 10999
rect 15577 10965 15611 10999
rect 16037 10965 16071 10999
rect 2789 10761 2823 10795
rect 3709 10761 3743 10795
rect 4077 10761 4111 10795
rect 7941 10761 7975 10795
rect 9413 10761 9447 10795
rect 10793 10761 10827 10795
rect 11713 10761 11747 10795
rect 12081 10761 12115 10795
rect 13737 10761 13771 10795
rect 13829 10761 13863 10795
rect 1676 10693 1710 10727
rect 5825 10693 5859 10727
rect 5917 10693 5951 10727
rect 8300 10693 8334 10727
rect 12173 10693 12207 10727
rect 13369 10693 13403 10727
rect 14105 10693 14139 10727
rect 14197 10693 14231 10727
rect 1409 10625 1443 10659
rect 3617 10625 3651 10659
rect 4721 10625 4755 10659
rect 4997 10625 5031 10659
rect 5549 10625 5583 10659
rect 5697 10625 5731 10659
rect 6055 10625 6089 10659
rect 6561 10625 6595 10659
rect 6828 10625 6862 10659
rect 8033 10625 8067 10659
rect 9505 10625 9539 10659
rect 12541 10625 12575 10659
rect 13093 10625 13127 10659
rect 13241 10625 13275 10659
rect 13461 10625 13495 10659
rect 13558 10625 13592 10659
rect 13967 10625 14001 10659
rect 14325 10625 14359 10659
rect 14473 10625 14507 10659
rect 14749 10625 14783 10659
rect 16230 10625 16264 10659
rect 16497 10625 16531 10659
rect 17049 10625 17083 10659
rect 17693 10625 17727 10659
rect 3433 10557 3467 10591
rect 12265 10557 12299 10591
rect 13001 10557 13035 10591
rect 17141 10557 17175 10591
rect 17325 10557 17359 10591
rect 5457 10489 5491 10523
rect 15117 10489 15151 10523
rect 17509 10489 17543 10523
rect 4169 10421 4203 10455
rect 5273 10421 5307 10455
rect 6193 10421 6227 10455
rect 12633 10421 12667 10455
rect 14565 10421 14599 10455
rect 16681 10421 16715 10455
rect 1501 10217 1535 10251
rect 2237 10217 2271 10251
rect 7297 10217 7331 10251
rect 9965 10217 9999 10251
rect 12265 10217 12299 10251
rect 12817 10217 12851 10251
rect 13921 10217 13955 10251
rect 14841 10217 14875 10251
rect 16037 10217 16071 10251
rect 17509 10217 17543 10251
rect 2789 10081 2823 10115
rect 10609 10081 10643 10115
rect 11345 10081 11379 10115
rect 14289 10081 14323 10115
rect 16865 10081 16899 10115
rect 1685 10013 1719 10047
rect 2053 10013 2087 10047
rect 2605 10013 2639 10047
rect 7481 10013 7515 10047
rect 7573 10013 7607 10047
rect 10333 10013 10367 10047
rect 12155 10013 12189 10047
rect 13277 10013 13311 10047
rect 13461 10013 13495 10047
rect 13737 10013 13771 10047
rect 15485 10013 15519 10047
rect 15853 10013 15887 10047
rect 11621 9945 11655 9979
rect 11989 9945 12023 9979
rect 12725 9945 12759 9979
rect 14381 9945 14415 9979
rect 14933 9945 14967 9979
rect 1869 9877 1903 9911
rect 2697 9877 2731 9911
rect 7757 9877 7791 9911
rect 10425 9877 10459 9911
rect 10793 9877 10827 9911
rect 14473 9877 14507 9911
rect 13277 9673 13311 9707
rect 13461 9673 13495 9707
rect 6377 9605 6411 9639
rect 10358 9605 10392 9639
rect 13001 9605 13035 9639
rect 14574 9605 14608 9639
rect 2237 9537 2271 9571
rect 2697 9537 2731 9571
rect 3781 9537 3815 9571
rect 6561 9537 6595 9571
rect 7941 9537 7975 9571
rect 8953 9537 8987 9571
rect 9045 9537 9079 9571
rect 10241 9537 10275 9571
rect 10793 9537 10827 9571
rect 11621 9537 11655 9571
rect 12265 9537 12299 9571
rect 1685 9469 1719 9503
rect 2789 9469 2823 9503
rect 2881 9469 2915 9503
rect 3525 9469 3559 9503
rect 5549 9469 5583 9503
rect 6837 9469 6871 9503
rect 7021 9469 7055 9503
rect 8217 9469 8251 9503
rect 8493 9469 8527 9503
rect 9413 9469 9447 9503
rect 9505 9469 9539 9503
rect 9873 9469 9907 9503
rect 10149 9469 10183 9503
rect 11897 9469 11931 9503
rect 14841 9469 14875 9503
rect 15945 9469 15979 9503
rect 17233 9469 17267 9503
rect 4905 9401 4939 9435
rect 8125 9401 8159 9435
rect 10517 9401 10551 9435
rect 16681 9401 16715 9435
rect 2329 9333 2363 9367
rect 4997 9333 5031 9367
rect 6745 9333 6779 9367
rect 7665 9333 7699 9367
rect 7757 9333 7791 9367
rect 10885 9333 10919 9367
rect 12081 9333 12115 9367
rect 16497 9333 16531 9367
rect 6561 9129 6595 9163
rect 6653 9129 6687 9163
rect 8677 9129 8711 9163
rect 10793 9129 10827 9163
rect 11437 9129 11471 9163
rect 14289 9129 14323 9163
rect 16405 9129 16439 9163
rect 3525 9061 3559 9095
rect 13093 9061 13127 9095
rect 14933 9061 14967 9095
rect 4537 8993 4571 9027
rect 5365 8993 5399 9027
rect 5641 8993 5675 9027
rect 5917 8993 5951 9027
rect 8493 8993 8527 9027
rect 9045 8993 9079 9027
rect 10517 8993 10551 9027
rect 10885 8993 10919 9027
rect 13829 8993 13863 9027
rect 16589 8993 16623 9027
rect 1777 8925 1811 8959
rect 1869 8925 1903 8959
rect 2145 8925 2179 8959
rect 4261 8925 4295 8959
rect 4721 8925 4755 8959
rect 4905 8925 4939 8959
rect 5779 8925 5813 8959
rect 7766 8925 7800 8959
rect 8033 8925 8067 8959
rect 8309 8925 8343 8959
rect 9505 8925 9539 8959
rect 10057 8925 10091 8959
rect 10149 8925 10183 8959
rect 11253 8925 11287 8959
rect 11713 8925 11747 8959
rect 14565 8925 14599 8959
rect 14749 8925 14783 8959
rect 15025 8925 15059 8959
rect 16865 8925 16899 8959
rect 17325 8925 17359 8959
rect 2390 8857 2424 8891
rect 4353 8857 4387 8891
rect 8769 8857 8803 8891
rect 9137 8857 9171 8891
rect 9597 8857 9631 8891
rect 10425 8857 10459 8891
rect 10634 8857 10668 8891
rect 11980 8857 12014 8891
rect 15270 8857 15304 8891
rect 1593 8789 1627 8823
rect 2053 8789 2087 8823
rect 3893 8789 3927 8823
rect 8125 8789 8159 8823
rect 11069 8789 11103 8823
rect 11161 8789 11195 8823
rect 13185 8789 13219 8823
rect 14105 8789 14139 8823
rect 16773 8789 16807 8823
rect 17233 8789 17267 8823
rect 17509 8789 17543 8823
rect 2973 8585 3007 8619
rect 3433 8585 3467 8619
rect 3985 8585 4019 8619
rect 6193 8585 6227 8619
rect 7297 8585 7331 8619
rect 8401 8585 8435 8619
rect 10517 8585 10551 8619
rect 11989 8585 12023 8619
rect 12357 8585 12391 8619
rect 13553 8585 13587 8619
rect 15209 8585 15243 8619
rect 15669 8585 15703 8619
rect 8125 8517 8159 8551
rect 8769 8517 8803 8551
rect 9229 8517 9263 8551
rect 10793 8517 10827 8551
rect 12449 8517 12483 8551
rect 1409 8449 1443 8483
rect 1676 8449 1710 8483
rect 3341 8449 3375 8483
rect 4169 8449 4203 8483
rect 4353 8449 4387 8483
rect 5390 8449 5424 8483
rect 7205 8449 7239 8483
rect 9137 8449 9171 8483
rect 9689 8449 9723 8483
rect 9873 8449 9907 8483
rect 10358 8449 10392 8483
rect 13277 8449 13311 8483
rect 14105 8449 14139 8483
rect 14381 8449 14415 8483
rect 14565 8449 14599 8483
rect 15577 8449 15611 8483
rect 16865 8449 16899 8483
rect 17233 8449 17267 8483
rect 3617 8381 3651 8415
rect 4537 8381 4571 8415
rect 5273 8381 5307 8415
rect 5549 8381 5583 8415
rect 7021 8381 7055 8415
rect 8677 8381 8711 8415
rect 10149 8381 10183 8415
rect 10241 8381 10275 8415
rect 12541 8381 12575 8415
rect 15761 8381 15795 8415
rect 16313 8381 16347 8415
rect 16957 8381 16991 8415
rect 2789 8313 2823 8347
rect 4997 8313 5031 8347
rect 7665 8313 7699 8347
rect 16681 8313 16715 8347
rect 10885 8245 10919 8279
rect 13921 8245 13955 8279
rect 3801 8041 3835 8075
rect 10793 8041 10827 8075
rect 12357 8041 12391 8075
rect 13001 8041 13035 8075
rect 16405 8041 16439 8075
rect 8217 7973 8251 8007
rect 4353 7905 4387 7939
rect 7573 7905 7607 7939
rect 5457 7837 5491 7871
rect 6929 7837 6963 7871
rect 7205 7837 7239 7871
rect 7389 7837 7423 7871
rect 7849 7837 7883 7871
rect 10701 7837 10735 7871
rect 12541 7837 12575 7871
rect 12730 7847 12764 7881
rect 13461 7837 13495 7871
rect 13737 7837 13771 7871
rect 13921 7837 13955 7871
rect 14381 7837 14415 7871
rect 17785 7837 17819 7871
rect 4813 7769 4847 7803
rect 13277 7769 13311 7803
rect 17518 7769 17552 7803
rect 5273 7701 5307 7735
rect 6745 7701 6779 7735
rect 7757 7701 7791 7735
rect 11161 7701 11195 7735
rect 13185 7701 13219 7735
rect 15669 7701 15703 7735
rect 7297 7497 7331 7531
rect 13829 7497 13863 7531
rect 14197 7497 14231 7531
rect 3341 7429 3375 7463
rect 6193 7429 6227 7463
rect 7389 7429 7423 7463
rect 10701 7429 10735 7463
rect 13461 7429 13495 7463
rect 3249 7361 3283 7395
rect 3709 7361 3743 7395
rect 4445 7361 4479 7395
rect 9485 7361 9519 7395
rect 11713 7361 11747 7395
rect 11989 7361 12023 7395
rect 12173 7361 12207 7395
rect 12357 7361 12391 7395
rect 12505 7361 12539 7395
rect 12633 7361 12667 7395
rect 12725 7361 12759 7395
rect 12822 7361 12856 7395
rect 13093 7361 13127 7395
rect 13241 7361 13275 7395
rect 13369 7361 13403 7395
rect 13599 7361 13633 7395
rect 16241 7361 16275 7395
rect 16497 7361 16531 7395
rect 17785 7361 17819 7395
rect 3433 7293 3467 7327
rect 4261 7293 4295 7327
rect 6745 7293 6779 7327
rect 9229 7293 9263 7327
rect 11253 7293 11287 7327
rect 14289 7293 14323 7327
rect 14473 7293 14507 7327
rect 14657 7293 14691 7327
rect 17509 7293 17543 7327
rect 15117 7225 15151 7259
rect 2881 7157 2915 7191
rect 8677 7157 8711 7191
rect 10609 7157 10643 7191
rect 11529 7157 11563 7191
rect 13001 7157 13035 7191
rect 13737 7157 13771 7191
rect 5549 6953 5583 6987
rect 7389 6953 7423 6987
rect 10241 6953 10275 6987
rect 14105 6953 14139 6987
rect 15025 6953 15059 6987
rect 9689 6817 9723 6851
rect 14657 6817 14691 6851
rect 15485 6817 15519 6851
rect 16405 6817 16439 6851
rect 2053 6749 2087 6783
rect 4169 6749 4203 6783
rect 4436 6749 4470 6783
rect 5917 6749 5951 6783
rect 6065 6749 6099 6783
rect 6423 6749 6457 6783
rect 6653 6749 6687 6783
rect 6837 6749 6871 6783
rect 7113 6749 7147 6783
rect 7297 6749 7331 6783
rect 8769 6749 8803 6783
rect 9505 6749 9539 6783
rect 9965 6749 9999 6783
rect 10517 6749 10551 6783
rect 10610 6749 10644 6783
rect 11021 6749 11055 6783
rect 11253 6749 11287 6783
rect 11437 6749 11471 6783
rect 11713 6749 11747 6783
rect 11897 6749 11931 6783
rect 13921 6749 13955 6783
rect 14473 6749 14507 6783
rect 15209 6749 15243 6783
rect 2320 6681 2354 6715
rect 6193 6681 6227 6715
rect 6285 6681 6319 6715
rect 8502 6681 8536 6715
rect 10793 6681 10827 6715
rect 10885 6681 10919 6715
rect 14565 6681 14599 6715
rect 16672 6681 16706 6715
rect 3433 6613 3467 6647
rect 6561 6613 6595 6647
rect 9137 6613 9171 6647
rect 9597 6613 9631 6647
rect 10425 6613 10459 6647
rect 11161 6613 11195 6647
rect 12633 6613 12667 6647
rect 15669 6613 15703 6647
rect 15761 6613 15795 6647
rect 16129 6613 16163 6647
rect 17785 6613 17819 6647
rect 2513 6409 2547 6443
rect 3341 6409 3375 6443
rect 4169 6409 4203 6443
rect 4537 6409 4571 6443
rect 4997 6409 5031 6443
rect 5457 6409 5491 6443
rect 9137 6409 9171 6443
rect 11621 6409 11655 6443
rect 15669 6409 15703 6443
rect 16497 6409 16531 6443
rect 16681 6409 16715 6443
rect 6745 6341 6779 6375
rect 11069 6341 11103 6375
rect 12081 6341 12115 6375
rect 16037 6341 16071 6375
rect 2697 6273 2731 6307
rect 5089 6273 5123 6307
rect 5549 6273 5583 6307
rect 6556 6273 6590 6307
rect 6653 6273 6687 6307
rect 6900 6273 6934 6307
rect 7021 6273 7055 6307
rect 7573 6273 7607 6307
rect 8033 6273 8067 6307
rect 8953 6273 8987 6307
rect 10701 6273 10735 6307
rect 10794 6273 10828 6307
rect 10977 6273 11011 6307
rect 11166 6273 11200 6307
rect 11989 6273 12023 6307
rect 12633 6273 12667 6307
rect 15025 6273 15059 6307
rect 16129 6273 16163 6307
rect 16865 6273 16899 6307
rect 17785 6273 17819 6307
rect 3157 6205 3191 6239
rect 3249 6205 3283 6239
rect 3985 6205 4019 6239
rect 4077 6205 4111 6239
rect 4813 6205 4847 6239
rect 6193 6205 6227 6239
rect 7665 6205 7699 6239
rect 12265 6205 12299 6239
rect 15853 6205 15887 6239
rect 17509 6205 17543 6239
rect 3709 6137 3743 6171
rect 7113 6137 7147 6171
rect 6377 6069 6411 6103
rect 7297 6069 7331 6103
rect 8217 6069 8251 6103
rect 11345 6069 11379 6103
rect 3617 5865 3651 5899
rect 5825 5865 5859 5899
rect 6009 5865 6043 5899
rect 12817 5865 12851 5899
rect 14933 5865 14967 5899
rect 3801 5797 3835 5831
rect 8769 5797 8803 5831
rect 16405 5797 16439 5831
rect 4445 5729 4479 5763
rect 5181 5729 5215 5763
rect 6561 5729 6595 5763
rect 7113 5729 7147 5763
rect 9505 5729 9539 5763
rect 10701 5729 10735 5763
rect 10793 5729 10827 5763
rect 11345 5729 11379 5763
rect 13277 5729 13311 5763
rect 13369 5729 13403 5763
rect 14381 5729 14415 5763
rect 15761 5729 15795 5763
rect 15945 5729 15979 5763
rect 17785 5729 17819 5763
rect 3433 5661 3467 5695
rect 5549 5661 5583 5695
rect 6285 5661 6319 5695
rect 6469 5661 6503 5695
rect 6837 5661 6871 5695
rect 7021 5661 7055 5695
rect 7389 5661 7423 5695
rect 10977 5661 11011 5695
rect 11253 5661 11287 5695
rect 11529 5661 11563 5695
rect 12265 5661 12299 5695
rect 13185 5661 13219 5695
rect 14565 5661 14599 5695
rect 15393 5661 15427 5695
rect 16497 5661 16531 5695
rect 17509 5661 17543 5695
rect 4169 5593 4203 5627
rect 4629 5593 4663 5627
rect 7656 5593 7690 5627
rect 11161 5593 11195 5627
rect 12541 5593 12575 5627
rect 15025 5593 15059 5627
rect 16037 5593 16071 5627
rect 4261 5525 4295 5559
rect 6101 5525 6135 5559
rect 6653 5525 6687 5559
rect 8953 5525 8987 5559
rect 11713 5525 11747 5559
rect 15209 5525 15243 5559
rect 16681 5525 16715 5559
rect 3985 5321 4019 5355
rect 8217 5321 8251 5355
rect 8769 5321 8803 5355
rect 11069 5321 11103 5355
rect 16129 5321 16163 5355
rect 4344 5253 4378 5287
rect 15016 5253 15050 5287
rect 2605 5185 2639 5219
rect 2872 5185 2906 5219
rect 6193 5185 6227 5219
rect 7297 5185 7331 5219
rect 7573 5185 7607 5219
rect 11713 5185 11747 5219
rect 13737 5185 13771 5219
rect 13854 5185 13888 5219
rect 17417 5185 17451 5219
rect 4077 5117 4111 5151
rect 6377 5117 6411 5151
rect 6561 5117 6595 5151
rect 7414 5117 7448 5151
rect 8861 5117 8895 5151
rect 9045 5117 9079 5151
rect 9229 5117 9263 5151
rect 9413 5117 9447 5151
rect 10149 5117 10183 5151
rect 10266 5117 10300 5151
rect 10425 5117 10459 5151
rect 12817 5117 12851 5151
rect 13001 5117 13035 5151
rect 14013 5117 14047 5151
rect 14749 5117 14783 5151
rect 17325 5117 17359 5151
rect 5457 5049 5491 5083
rect 7021 5049 7055 5083
rect 9873 5049 9907 5083
rect 13461 5049 13495 5083
rect 5549 4981 5583 5015
rect 8401 4981 8435 5015
rect 11529 4981 11563 5015
rect 14657 4981 14691 5015
rect 16681 4981 16715 5015
rect 17601 4981 17635 5015
rect 2973 4777 3007 4811
rect 4537 4777 4571 4811
rect 5641 4777 5675 4811
rect 8125 4777 8159 4811
rect 11069 4777 11103 4811
rect 13553 4777 13587 4811
rect 13921 4777 13955 4811
rect 15025 4777 15059 4811
rect 17693 4777 17727 4811
rect 6837 4709 6871 4743
rect 12633 4709 12667 4743
rect 14933 4709 14967 4743
rect 4997 4641 5031 4675
rect 5181 4641 5215 4675
rect 6275 4641 6309 4675
rect 6542 4641 6576 4675
rect 7481 4641 7515 4675
rect 9413 4641 9447 4675
rect 9873 4641 9907 4675
rect 10266 4641 10300 4675
rect 10425 4641 10459 4675
rect 13369 4641 13403 4675
rect 15669 4641 15703 4675
rect 3157 4573 3191 4607
rect 4905 4573 4939 4607
rect 6423 4573 6457 4607
rect 7297 4573 7331 4607
rect 8309 4573 8343 4607
rect 9229 4573 9263 4607
rect 10149 4573 10183 4607
rect 11253 4573 11287 4607
rect 13461 4573 13495 4607
rect 13737 4573 13771 4607
rect 14473 4573 14507 4607
rect 14565 4573 14599 4607
rect 14749 4573 14783 4607
rect 15393 4573 15427 4607
rect 17325 4573 17359 4607
rect 17509 4573 17543 4607
rect 11498 4505 11532 4539
rect 17058 4505 17092 4539
rect 12725 4437 12759 4471
rect 15485 4437 15519 4471
rect 15945 4437 15979 4471
rect 11713 4233 11747 4267
rect 12081 4233 12115 4267
rect 14657 4233 14691 4267
rect 6745 4165 6779 4199
rect 7205 4165 7239 4199
rect 15577 4165 15611 4199
rect 6837 4097 6871 4131
rect 7757 4097 7791 4131
rect 10517 4097 10551 4131
rect 12725 4097 12759 4131
rect 12817 4097 12851 4131
rect 13737 4097 13771 4131
rect 13854 4097 13888 4131
rect 14013 4097 14047 4131
rect 15209 4097 15243 4131
rect 15853 4097 15887 4131
rect 16957 4097 16991 4131
rect 17509 4097 17543 4131
rect 5825 4029 5859 4063
rect 7021 4029 7055 4063
rect 8769 4029 8803 4063
rect 12173 4029 12207 4063
rect 12265 4029 12299 4063
rect 13001 4029 13035 4063
rect 13461 4029 13495 4063
rect 16405 4029 16439 4063
rect 5273 3893 5307 3927
rect 6377 3893 6411 3927
rect 8125 3893 8159 3927
rect 11161 3893 11195 3927
rect 12541 3893 12575 3927
rect 6745 3689 6779 3723
rect 4537 3621 4571 3655
rect 8769 3621 8803 3655
rect 10609 3621 10643 3655
rect 13001 3621 13035 3655
rect 14841 3621 14875 3655
rect 4997 3553 5031 3587
rect 5181 3553 5215 3587
rect 7113 3553 7147 3587
rect 8217 3553 8251 3587
rect 10149 3553 10183 3587
rect 11161 3553 11195 3587
rect 12357 3553 12391 3587
rect 12541 3553 12575 3587
rect 13737 3553 13771 3587
rect 15301 3553 15335 3587
rect 15393 3553 15427 3587
rect 4445 3485 4479 3519
rect 4905 3485 4939 3519
rect 5365 3485 5399 3519
rect 7297 3485 7331 3519
rect 8401 3485 8435 3519
rect 9137 3485 9171 3519
rect 9413 3485 9447 3519
rect 10977 3485 11011 3519
rect 11989 3485 12023 3519
rect 14105 3485 14139 3519
rect 14565 3485 14599 3519
rect 16221 3485 16255 3519
rect 5632 3417 5666 3451
rect 8309 3417 8343 3451
rect 9873 3417 9907 3451
rect 11437 3417 11471 3451
rect 12633 3417 12667 3451
rect 13093 3417 13127 3451
rect 15209 3417 15243 3451
rect 15669 3417 15703 3451
rect 17693 3417 17727 3451
rect 4261 3349 4295 3383
rect 7205 3349 7239 3383
rect 7665 3349 7699 3383
rect 8953 3349 8987 3383
rect 9229 3349 9263 3383
rect 9505 3349 9539 3383
rect 9965 3349 9999 3383
rect 11069 3349 11103 3383
rect 14289 3349 14323 3383
rect 14749 3349 14783 3383
rect 17601 3349 17635 3383
rect 5549 3145 5583 3179
rect 5641 3145 5675 3179
rect 6377 3145 6411 3179
rect 9229 3145 9263 3179
rect 9873 3145 9907 3179
rect 9965 3145 9999 3179
rect 13185 3145 13219 3179
rect 16037 3145 16071 3179
rect 4414 3077 4448 3111
rect 8116 3077 8150 3111
rect 11078 3077 11112 3111
rect 14902 3077 14936 3111
rect 4169 3009 4203 3043
rect 5825 3009 5859 3043
rect 7501 3009 7535 3043
rect 7757 3009 7791 3043
rect 7849 3009 7883 3043
rect 9413 3009 9447 3043
rect 9689 3009 9723 3043
rect 11345 3009 11379 3043
rect 11713 3009 11747 3043
rect 11980 3009 12014 3043
rect 14298 3009 14332 3043
rect 14565 3009 14599 3043
rect 14657 3009 14691 3043
rect 9505 2805 9539 2839
rect 13093 2805 13127 2839
rect 7573 2601 7607 2635
rect 7665 2601 7699 2635
rect 10425 2601 10459 2635
rect 14105 2601 14139 2635
rect 4261 2533 4295 2567
rect 13001 2533 13035 2567
rect 13461 2533 13495 2567
rect 6929 2465 6963 2499
rect 9045 2465 9079 2499
rect 10793 2465 10827 2499
rect 11805 2465 11839 2499
rect 14565 2465 14599 2499
rect 14657 2465 14691 2499
rect 5917 2397 5951 2431
rect 6561 2397 6595 2431
rect 7849 2397 7883 2431
rect 8493 2397 8527 2431
rect 8769 2397 8803 2431
rect 9312 2397 9346 2431
rect 10517 2397 10551 2431
rect 11529 2397 11563 2431
rect 12449 2397 12483 2431
rect 12817 2397 12851 2431
rect 15485 2397 15519 2431
rect 4077 2329 4111 2363
rect 13277 2329 13311 2363
rect 14473 2329 14507 2363
rect 14933 2329 14967 2363
rect 6101 2261 6135 2295
rect 6745 2261 6779 2295
rect 12633 2261 12667 2295
<< metal1 >>
rect 1104 19066 18124 19088
rect 1104 19014 3077 19066
rect 3129 19014 3141 19066
rect 3193 19014 3205 19066
rect 3257 19014 3269 19066
rect 3321 19014 3333 19066
rect 3385 19014 7332 19066
rect 7384 19014 7396 19066
rect 7448 19014 7460 19066
rect 7512 19014 7524 19066
rect 7576 19014 7588 19066
rect 7640 19014 11587 19066
rect 11639 19014 11651 19066
rect 11703 19014 11715 19066
rect 11767 19014 11779 19066
rect 11831 19014 11843 19066
rect 11895 19014 15842 19066
rect 15894 19014 15906 19066
rect 15958 19014 15970 19066
rect 16022 19014 16034 19066
rect 16086 19014 16098 19066
rect 16150 19014 18124 19066
rect 1104 18992 18124 19014
rect 10045 18955 10103 18961
rect 10045 18921 10057 18955
rect 10091 18952 10103 18955
rect 10318 18952 10324 18964
rect 10091 18924 10324 18952
rect 10091 18921 10103 18924
rect 10045 18915 10103 18921
rect 10318 18912 10324 18924
rect 10376 18912 10382 18964
rect 12618 18912 12624 18964
rect 12676 18912 12682 18964
rect 7098 18708 7104 18760
rect 7156 18708 7162 18760
rect 7469 18751 7527 18757
rect 7469 18717 7481 18751
rect 7515 18748 7527 18751
rect 7834 18748 7840 18760
rect 7515 18720 7840 18748
rect 7515 18717 7527 18720
rect 7469 18711 7527 18717
rect 7834 18708 7840 18720
rect 7892 18708 7898 18760
rect 8389 18751 8447 18757
rect 8389 18717 8401 18751
rect 8435 18748 8447 18751
rect 8570 18748 8576 18760
rect 8435 18720 8576 18748
rect 8435 18717 8447 18720
rect 8389 18711 8447 18717
rect 8570 18708 8576 18720
rect 8628 18708 8634 18760
rect 8665 18751 8723 18757
rect 8665 18717 8677 18751
rect 8711 18748 8723 18751
rect 9030 18748 9036 18760
rect 8711 18720 9036 18748
rect 8711 18717 8723 18720
rect 8665 18711 8723 18717
rect 9030 18708 9036 18720
rect 9088 18708 9094 18760
rect 9306 18708 9312 18760
rect 9364 18748 9370 18760
rect 9493 18751 9551 18757
rect 9493 18748 9505 18751
rect 9364 18720 9505 18748
rect 9364 18708 9370 18720
rect 9493 18717 9505 18720
rect 9539 18717 9551 18751
rect 9493 18711 9551 18717
rect 10594 18708 10600 18760
rect 10652 18748 10658 18760
rect 10781 18751 10839 18757
rect 10781 18748 10793 18751
rect 10652 18720 10793 18748
rect 10652 18708 10658 18720
rect 10781 18717 10793 18720
rect 10827 18717 10839 18751
rect 10781 18711 10839 18717
rect 11146 18708 11152 18760
rect 11204 18708 11210 18760
rect 12161 18751 12219 18757
rect 12161 18717 12173 18751
rect 12207 18748 12219 18751
rect 12618 18748 12624 18760
rect 12207 18720 12624 18748
rect 12207 18717 12219 18720
rect 12161 18711 12219 18717
rect 12618 18708 12624 18720
rect 12676 18708 12682 18760
rect 13078 18708 13084 18760
rect 13136 18748 13142 18760
rect 13449 18751 13507 18757
rect 13449 18748 13461 18751
rect 13136 18720 13461 18748
rect 13136 18708 13142 18720
rect 13449 18717 13461 18720
rect 13495 18717 13507 18751
rect 13449 18711 13507 18717
rect 13814 18708 13820 18760
rect 13872 18708 13878 18760
rect 8478 18640 8484 18692
rect 8536 18640 8542 18692
rect 9766 18640 9772 18692
rect 9824 18640 9830 18692
rect 12713 18683 12771 18689
rect 12713 18649 12725 18683
rect 12759 18680 12771 18683
rect 14090 18680 14096 18692
rect 12759 18652 14096 18680
rect 12759 18649 12771 18652
rect 12713 18643 12771 18649
rect 14090 18640 14096 18652
rect 14148 18640 14154 18692
rect 6730 18572 6736 18624
rect 6788 18612 6794 18624
rect 6917 18615 6975 18621
rect 6917 18612 6929 18615
rect 6788 18584 6929 18612
rect 6788 18572 6794 18584
rect 6917 18581 6929 18584
rect 6963 18581 6975 18615
rect 6917 18575 6975 18581
rect 7650 18572 7656 18624
rect 7708 18572 7714 18624
rect 7742 18572 7748 18624
rect 7800 18572 7806 18624
rect 8938 18572 8944 18624
rect 8996 18572 9002 18624
rect 9858 18572 9864 18624
rect 9916 18612 9922 18624
rect 10229 18615 10287 18621
rect 10229 18612 10241 18615
rect 9916 18584 10241 18612
rect 9916 18572 9922 18584
rect 10229 18581 10241 18584
rect 10275 18581 10287 18615
rect 10229 18575 10287 18581
rect 11330 18572 11336 18624
rect 11388 18572 11394 18624
rect 11422 18572 11428 18624
rect 11480 18612 11486 18624
rect 11517 18615 11575 18621
rect 11517 18612 11529 18615
rect 11480 18584 11529 18612
rect 11480 18572 11486 18584
rect 11517 18581 11529 18584
rect 11563 18581 11575 18615
rect 11517 18575 11575 18581
rect 12894 18572 12900 18624
rect 12952 18572 12958 18624
rect 13630 18572 13636 18624
rect 13688 18572 13694 18624
rect 1104 18522 18124 18544
rect 1104 18470 3737 18522
rect 3789 18470 3801 18522
rect 3853 18470 3865 18522
rect 3917 18470 3929 18522
rect 3981 18470 3993 18522
rect 4045 18470 7992 18522
rect 8044 18470 8056 18522
rect 8108 18470 8120 18522
rect 8172 18470 8184 18522
rect 8236 18470 8248 18522
rect 8300 18470 12247 18522
rect 12299 18470 12311 18522
rect 12363 18470 12375 18522
rect 12427 18470 12439 18522
rect 12491 18470 12503 18522
rect 12555 18470 16502 18522
rect 16554 18470 16566 18522
rect 16618 18470 16630 18522
rect 16682 18470 16694 18522
rect 16746 18470 16758 18522
rect 16810 18470 18124 18522
rect 1104 18448 18124 18470
rect 7650 18368 7656 18420
rect 7708 18408 7714 18420
rect 7708 18380 7972 18408
rect 7708 18368 7714 18380
rect 7944 18340 7972 18380
rect 9306 18368 9312 18420
rect 9364 18368 9370 18420
rect 9493 18411 9551 18417
rect 9493 18377 9505 18411
rect 9539 18408 9551 18411
rect 9674 18408 9680 18420
rect 9539 18380 9680 18408
rect 9539 18377 9551 18380
rect 9493 18371 9551 18377
rect 9674 18368 9680 18380
rect 9732 18368 9738 18420
rect 10502 18408 10508 18420
rect 9784 18380 10508 18408
rect 9784 18349 9812 18380
rect 10502 18368 10508 18380
rect 10560 18368 10566 18420
rect 11974 18368 11980 18420
rect 12032 18408 12038 18420
rect 13078 18408 13084 18420
rect 12032 18380 13084 18408
rect 12032 18368 12038 18380
rect 13078 18368 13084 18380
rect 13136 18368 13142 18420
rect 8174 18343 8232 18349
rect 8174 18340 8186 18343
rect 6472 18312 7788 18340
rect 7944 18312 8186 18340
rect 6472 18281 6500 18312
rect 6730 18281 6736 18284
rect 6457 18275 6515 18281
rect 6457 18241 6469 18275
rect 6503 18241 6515 18275
rect 6724 18272 6736 18281
rect 6691 18244 6736 18272
rect 6457 18235 6515 18241
rect 6724 18235 6736 18244
rect 6730 18232 6736 18235
rect 6788 18232 6794 18284
rect 7760 18216 7788 18312
rect 8174 18309 8186 18312
rect 8220 18309 8232 18343
rect 8174 18303 8232 18309
rect 9769 18343 9827 18349
rect 9769 18309 9781 18343
rect 9815 18309 9827 18343
rect 11054 18340 11060 18352
rect 9769 18303 9827 18309
rect 9968 18312 11060 18340
rect 9968 18281 9996 18312
rect 11054 18300 11060 18312
rect 11112 18340 11118 18352
rect 13532 18343 13590 18349
rect 11112 18312 12434 18340
rect 11112 18300 11118 18312
rect 9953 18275 10011 18281
rect 9953 18241 9965 18275
rect 9999 18241 10011 18275
rect 9953 18235 10011 18241
rect 10220 18275 10278 18281
rect 10220 18241 10232 18275
rect 10266 18272 10278 18275
rect 10686 18272 10692 18284
rect 10266 18244 10692 18272
rect 10266 18241 10278 18244
rect 10220 18235 10278 18241
rect 10686 18232 10692 18244
rect 10744 18232 10750 18284
rect 11716 18281 11744 18312
rect 11701 18275 11759 18281
rect 11701 18241 11713 18275
rect 11747 18241 11759 18275
rect 11957 18275 12015 18281
rect 11957 18272 11969 18275
rect 11701 18235 11759 18241
rect 11808 18244 11969 18272
rect 7742 18164 7748 18216
rect 7800 18204 7806 18216
rect 7929 18207 7987 18213
rect 7929 18204 7941 18207
rect 7800 18176 7941 18204
rect 7800 18164 7806 18176
rect 7929 18173 7941 18176
rect 7975 18173 7987 18207
rect 7929 18167 7987 18173
rect 11330 18164 11336 18216
rect 11388 18204 11394 18216
rect 11808 18204 11836 18244
rect 11957 18241 11969 18244
rect 12003 18241 12015 18275
rect 12406 18272 12434 18312
rect 13532 18309 13544 18343
rect 13578 18340 13590 18343
rect 13630 18340 13636 18352
rect 13578 18312 13636 18340
rect 13578 18309 13590 18312
rect 13532 18303 13590 18309
rect 13630 18300 13636 18312
rect 13688 18300 13694 18352
rect 13265 18275 13323 18281
rect 13265 18272 13277 18275
rect 12406 18244 13277 18272
rect 11957 18235 12015 18241
rect 13265 18241 13277 18244
rect 13311 18241 13323 18275
rect 13265 18235 13323 18241
rect 15654 18232 15660 18284
rect 15712 18232 15718 18284
rect 11388 18176 11836 18204
rect 15289 18207 15347 18213
rect 11388 18164 11394 18176
rect 15289 18173 15301 18207
rect 15335 18173 15347 18207
rect 15289 18167 15347 18173
rect 14645 18139 14703 18145
rect 14645 18105 14657 18139
rect 14691 18136 14703 18139
rect 15010 18136 15016 18148
rect 14691 18108 15016 18136
rect 14691 18105 14703 18108
rect 14645 18099 14703 18105
rect 15010 18096 15016 18108
rect 15068 18136 15074 18148
rect 15304 18136 15332 18167
rect 15068 18108 15332 18136
rect 15068 18096 15074 18108
rect 7837 18071 7895 18077
rect 7837 18037 7849 18071
rect 7883 18068 7895 18071
rect 8570 18068 8576 18080
rect 7883 18040 8576 18068
rect 7883 18037 7895 18040
rect 7837 18031 7895 18037
rect 8570 18028 8576 18040
rect 8628 18068 8634 18080
rect 9490 18068 9496 18080
rect 8628 18040 9496 18068
rect 8628 18028 8634 18040
rect 9490 18028 9496 18040
rect 9548 18028 9554 18080
rect 11333 18071 11391 18077
rect 11333 18037 11345 18071
rect 11379 18068 11391 18071
rect 12618 18068 12624 18080
rect 11379 18040 12624 18068
rect 11379 18037 11391 18040
rect 11333 18031 11391 18037
rect 12618 18028 12624 18040
rect 12676 18028 12682 18080
rect 14734 18028 14740 18080
rect 14792 18028 14798 18080
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 15473 18071 15531 18077
rect 15473 18068 15485 18071
rect 15436 18040 15485 18068
rect 15436 18028 15442 18040
rect 15473 18037 15485 18040
rect 15519 18037 15531 18071
rect 15473 18031 15531 18037
rect 1104 17978 18124 18000
rect 1104 17926 3077 17978
rect 3129 17926 3141 17978
rect 3193 17926 3205 17978
rect 3257 17926 3269 17978
rect 3321 17926 3333 17978
rect 3385 17926 7332 17978
rect 7384 17926 7396 17978
rect 7448 17926 7460 17978
rect 7512 17926 7524 17978
rect 7576 17926 7588 17978
rect 7640 17926 11587 17978
rect 11639 17926 11651 17978
rect 11703 17926 11715 17978
rect 11767 17926 11779 17978
rect 11831 17926 11843 17978
rect 11895 17926 15842 17978
rect 15894 17926 15906 17978
rect 15958 17926 15970 17978
rect 16022 17926 16034 17978
rect 16086 17926 16098 17978
rect 16150 17926 18124 17978
rect 1104 17904 18124 17926
rect 7098 17824 7104 17876
rect 7156 17864 7162 17876
rect 7193 17867 7251 17873
rect 7193 17864 7205 17867
rect 7156 17836 7205 17864
rect 7156 17824 7162 17836
rect 7193 17833 7205 17836
rect 7239 17833 7251 17867
rect 7193 17827 7251 17833
rect 7834 17824 7840 17876
rect 7892 17864 7898 17876
rect 8021 17867 8079 17873
rect 8021 17864 8033 17867
rect 7892 17836 8033 17864
rect 7892 17824 7898 17836
rect 8021 17833 8033 17836
rect 8067 17833 8079 17867
rect 8021 17827 8079 17833
rect 8680 17836 10088 17864
rect 8386 17796 8392 17808
rect 6932 17768 8392 17796
rect 5166 17688 5172 17740
rect 5224 17728 5230 17740
rect 6932 17737 6960 17768
rect 8386 17756 8392 17768
rect 8444 17756 8450 17808
rect 8680 17740 8708 17836
rect 10060 17796 10088 17836
rect 10134 17824 10140 17876
rect 10192 17864 10198 17876
rect 10505 17867 10563 17873
rect 10505 17864 10517 17867
rect 10192 17836 10517 17864
rect 10192 17824 10198 17836
rect 10505 17833 10517 17836
rect 10551 17864 10563 17867
rect 10594 17864 10600 17876
rect 10551 17836 10600 17864
rect 10551 17833 10563 17836
rect 10505 17827 10563 17833
rect 10594 17824 10600 17836
rect 10652 17824 10658 17876
rect 10686 17824 10692 17876
rect 10744 17824 10750 17876
rect 11146 17824 11152 17876
rect 11204 17864 11210 17876
rect 12161 17867 12219 17873
rect 12161 17864 12173 17867
rect 11204 17836 12173 17864
rect 11204 17824 11210 17836
rect 12161 17833 12173 17836
rect 12207 17833 12219 17867
rect 12161 17827 12219 17833
rect 13814 17824 13820 17876
rect 13872 17864 13878 17876
rect 13909 17867 13967 17873
rect 13909 17864 13921 17867
rect 13872 17836 13921 17864
rect 13872 17824 13878 17836
rect 13909 17833 13921 17836
rect 13955 17833 13967 17867
rect 13909 17827 13967 17833
rect 14277 17867 14335 17873
rect 14277 17833 14289 17867
rect 14323 17864 14335 17867
rect 14323 17836 16344 17864
rect 14323 17833 14335 17836
rect 14277 17827 14335 17833
rect 10060 17768 12020 17796
rect 6733 17731 6791 17737
rect 6733 17728 6745 17731
rect 5224 17700 6745 17728
rect 5224 17688 5230 17700
rect 6733 17697 6745 17700
rect 6779 17697 6791 17731
rect 6733 17691 6791 17697
rect 6917 17731 6975 17737
rect 6917 17697 6929 17731
rect 6963 17697 6975 17731
rect 7837 17731 7895 17737
rect 7837 17728 7849 17731
rect 6917 17691 6975 17697
rect 7024 17700 7849 17728
rect 4706 17620 4712 17672
rect 4764 17620 4770 17672
rect 5074 17620 5080 17672
rect 5132 17620 5138 17672
rect 5626 17620 5632 17672
rect 5684 17620 5690 17672
rect 7024 17660 7052 17700
rect 7837 17697 7849 17700
rect 7883 17728 7895 17731
rect 8570 17728 8576 17740
rect 7883 17700 8576 17728
rect 7883 17697 7895 17700
rect 7837 17691 7895 17697
rect 8570 17688 8576 17700
rect 8628 17688 8634 17740
rect 8662 17688 8668 17740
rect 8720 17688 8726 17740
rect 11514 17728 11520 17740
rect 10796 17700 11520 17728
rect 5736 17632 7052 17660
rect 7561 17663 7619 17669
rect 4430 17552 4436 17604
rect 4488 17592 4494 17604
rect 5736 17592 5764 17632
rect 7561 17629 7573 17663
rect 7607 17660 7619 17663
rect 7650 17660 7656 17672
rect 7607 17632 7656 17660
rect 7607 17629 7619 17632
rect 7561 17623 7619 17629
rect 7650 17620 7656 17632
rect 7708 17620 7714 17672
rect 7742 17620 7748 17672
rect 7800 17660 7806 17672
rect 9125 17663 9183 17669
rect 9125 17660 9137 17663
rect 7800 17632 9137 17660
rect 7800 17620 7806 17632
rect 9125 17629 9137 17632
rect 9171 17629 9183 17663
rect 9125 17623 9183 17629
rect 4488 17564 5764 17592
rect 6181 17595 6239 17601
rect 4488 17552 4494 17564
rect 6181 17561 6193 17595
rect 6227 17592 6239 17595
rect 6641 17595 6699 17601
rect 6641 17592 6653 17595
rect 6227 17564 6653 17592
rect 6227 17561 6239 17564
rect 6181 17555 6239 17561
rect 6641 17561 6653 17564
rect 6687 17561 6699 17595
rect 6641 17555 6699 17561
rect 8389 17595 8447 17601
rect 8389 17561 8401 17595
rect 8435 17592 8447 17595
rect 8938 17592 8944 17604
rect 8435 17564 8944 17592
rect 8435 17561 8447 17564
rect 8389 17555 8447 17561
rect 8938 17552 8944 17564
rect 8996 17552 9002 17604
rect 9392 17595 9450 17601
rect 9392 17561 9404 17595
rect 9438 17592 9450 17595
rect 10226 17592 10232 17604
rect 9438 17564 10232 17592
rect 9438 17561 9450 17564
rect 9392 17555 9450 17561
rect 10226 17552 10232 17564
rect 10284 17552 10290 17604
rect 4154 17484 4160 17536
rect 4212 17484 4218 17536
rect 4890 17484 4896 17536
rect 4948 17484 4954 17536
rect 5994 17484 6000 17536
rect 6052 17524 6058 17536
rect 6273 17527 6331 17533
rect 6273 17524 6285 17527
rect 6052 17496 6285 17524
rect 6052 17484 6058 17496
rect 6273 17493 6285 17496
rect 6319 17493 6331 17527
rect 6273 17487 6331 17493
rect 7653 17527 7711 17533
rect 7653 17493 7665 17527
rect 7699 17524 7711 17527
rect 8478 17524 8484 17536
rect 7699 17496 8484 17524
rect 7699 17493 7711 17496
rect 7653 17487 7711 17493
rect 8478 17484 8484 17496
rect 8536 17484 8542 17536
rect 8570 17484 8576 17536
rect 8628 17524 8634 17536
rect 10796 17524 10824 17700
rect 11514 17688 11520 17700
rect 11572 17688 11578 17740
rect 11992 17728 12020 17768
rect 12434 17756 12440 17808
rect 12492 17796 12498 17808
rect 12492 17768 13308 17796
rect 12492 17756 12498 17768
rect 12713 17731 12771 17737
rect 12713 17728 12725 17731
rect 11992 17700 12725 17728
rect 12713 17697 12725 17700
rect 12759 17728 12771 17731
rect 13170 17728 13176 17740
rect 12759 17700 13176 17728
rect 12759 17697 12771 17700
rect 12713 17691 12771 17697
rect 13170 17688 13176 17700
rect 13228 17688 13234 17740
rect 13280 17737 13308 17768
rect 13265 17731 13323 17737
rect 13265 17697 13277 17731
rect 13311 17697 13323 17731
rect 13265 17691 13323 17697
rect 16206 17688 16212 17740
rect 16264 17728 16270 17740
rect 16316 17737 16344 17836
rect 16301 17731 16359 17737
rect 16301 17728 16313 17731
rect 16264 17700 16313 17728
rect 16264 17688 16270 17700
rect 16301 17697 16313 17700
rect 16347 17697 16359 17731
rect 16301 17691 16359 17697
rect 10873 17663 10931 17669
rect 10873 17629 10885 17663
rect 10919 17660 10931 17663
rect 11333 17663 11391 17669
rect 10919 17632 11008 17660
rect 10919 17629 10931 17632
rect 10873 17623 10931 17629
rect 10980 17533 11008 17632
rect 11333 17629 11345 17663
rect 11379 17660 11391 17663
rect 11422 17660 11428 17672
rect 11379 17632 11428 17660
rect 11379 17629 11391 17632
rect 11333 17623 11391 17629
rect 11422 17620 11428 17632
rect 11480 17620 11486 17672
rect 11532 17660 11560 17688
rect 12434 17660 12440 17672
rect 11532 17632 12440 17660
rect 12434 17620 12440 17632
rect 12492 17620 12498 17672
rect 12529 17663 12587 17669
rect 12529 17629 12541 17663
rect 12575 17660 12587 17663
rect 12894 17660 12900 17672
rect 12575 17632 12900 17660
rect 12575 17629 12587 17632
rect 12529 17623 12587 17629
rect 12894 17620 12900 17632
rect 12952 17620 12958 17672
rect 14918 17660 14924 17672
rect 13464 17632 14924 17660
rect 13464 17592 13492 17632
rect 14918 17620 14924 17632
rect 14976 17620 14982 17672
rect 15378 17620 15384 17672
rect 15436 17669 15442 17672
rect 15436 17660 15448 17669
rect 15436 17632 15481 17660
rect 15436 17623 15448 17632
rect 15436 17620 15442 17623
rect 15562 17620 15568 17672
rect 15620 17660 15626 17672
rect 15657 17663 15715 17669
rect 15657 17660 15669 17663
rect 15620 17632 15669 17660
rect 15620 17620 15626 17632
rect 15657 17629 15669 17632
rect 15703 17629 15715 17663
rect 15657 17623 15715 17629
rect 12636 17564 13492 17592
rect 13541 17595 13599 17601
rect 8628 17496 10824 17524
rect 10965 17527 11023 17533
rect 8628 17484 8634 17496
rect 10965 17493 10977 17527
rect 11011 17493 11023 17527
rect 10965 17487 11023 17493
rect 11146 17484 11152 17536
rect 11204 17524 11210 17536
rect 12636 17533 12664 17564
rect 13541 17561 13553 17595
rect 13587 17592 13599 17595
rect 14734 17592 14740 17604
rect 13587 17564 14740 17592
rect 13587 17561 13599 17564
rect 13541 17555 13599 17561
rect 14734 17552 14740 17564
rect 14792 17552 14798 17604
rect 11425 17527 11483 17533
rect 11425 17524 11437 17527
rect 11204 17496 11437 17524
rect 11204 17484 11210 17496
rect 11425 17493 11437 17496
rect 11471 17524 11483 17527
rect 12621 17527 12679 17533
rect 12621 17524 12633 17527
rect 11471 17496 12633 17524
rect 11471 17493 11483 17496
rect 11425 17487 11483 17493
rect 12621 17493 12633 17496
rect 12667 17493 12679 17527
rect 12621 17487 12679 17493
rect 13449 17527 13507 17533
rect 13449 17493 13461 17527
rect 13495 17524 13507 17527
rect 14458 17524 14464 17536
rect 13495 17496 14464 17524
rect 13495 17493 13507 17496
rect 13449 17487 13507 17493
rect 14458 17484 14464 17496
rect 14516 17484 14522 17536
rect 14550 17484 14556 17536
rect 14608 17524 14614 17536
rect 15749 17527 15807 17533
rect 15749 17524 15761 17527
rect 14608 17496 15761 17524
rect 14608 17484 14614 17496
rect 15749 17493 15761 17496
rect 15795 17493 15807 17527
rect 15749 17487 15807 17493
rect 1104 17434 18124 17456
rect 1104 17382 3737 17434
rect 3789 17382 3801 17434
rect 3853 17382 3865 17434
rect 3917 17382 3929 17434
rect 3981 17382 3993 17434
rect 4045 17382 7992 17434
rect 8044 17382 8056 17434
rect 8108 17382 8120 17434
rect 8172 17382 8184 17434
rect 8236 17382 8248 17434
rect 8300 17382 12247 17434
rect 12299 17382 12311 17434
rect 12363 17382 12375 17434
rect 12427 17382 12439 17434
rect 12491 17382 12503 17434
rect 12555 17382 16502 17434
rect 16554 17382 16566 17434
rect 16618 17382 16630 17434
rect 16682 17382 16694 17434
rect 16746 17382 16758 17434
rect 16810 17382 18124 17434
rect 1104 17360 18124 17382
rect 3973 17323 4031 17329
rect 3973 17289 3985 17323
rect 4019 17320 4031 17323
rect 4706 17320 4712 17332
rect 4019 17292 4712 17320
rect 4019 17289 4031 17292
rect 3973 17283 4031 17289
rect 4706 17280 4712 17292
rect 4764 17320 4770 17332
rect 5258 17320 5264 17332
rect 4764 17292 5264 17320
rect 4764 17280 4770 17292
rect 5258 17280 5264 17292
rect 5316 17280 5322 17332
rect 6181 17323 6239 17329
rect 6181 17289 6193 17323
rect 6227 17289 6239 17323
rect 6181 17283 6239 17289
rect 9769 17323 9827 17329
rect 9769 17289 9781 17323
rect 9815 17320 9827 17323
rect 9858 17320 9864 17332
rect 9815 17292 9864 17320
rect 9815 17289 9827 17292
rect 9769 17283 9827 17289
rect 4516 17255 4574 17261
rect 4516 17221 4528 17255
rect 4562 17252 4574 17255
rect 4890 17252 4896 17264
rect 4562 17224 4896 17252
rect 4562 17221 4574 17224
rect 4516 17215 4574 17221
rect 4890 17212 4896 17224
rect 4948 17212 4954 17264
rect 2866 17193 2872 17196
rect 2860 17147 2872 17193
rect 2866 17144 2872 17147
rect 2924 17144 2930 17196
rect 5994 17144 6000 17196
rect 6052 17144 6058 17196
rect 6196 17184 6224 17283
rect 9858 17280 9864 17292
rect 9916 17280 9922 17332
rect 10226 17280 10232 17332
rect 10284 17280 10290 17332
rect 14458 17280 14464 17332
rect 14516 17280 14522 17332
rect 14550 17280 14556 17332
rect 14608 17280 14614 17332
rect 14921 17323 14979 17329
rect 14921 17289 14933 17323
rect 14967 17320 14979 17323
rect 15654 17320 15660 17332
rect 14967 17292 15660 17320
rect 14967 17289 14979 17292
rect 14921 17283 14979 17289
rect 15654 17280 15660 17292
rect 15712 17280 15718 17332
rect 10870 17252 10876 17264
rect 10060 17224 10876 17252
rect 7478 17187 7536 17193
rect 7478 17184 7490 17187
rect 6196 17156 7490 17184
rect 7478 17153 7490 17156
rect 7524 17153 7536 17187
rect 7478 17147 7536 17153
rect 7834 17144 7840 17196
rect 7892 17184 7898 17196
rect 8478 17184 8484 17196
rect 7892 17156 8484 17184
rect 7892 17144 7898 17156
rect 8478 17144 8484 17156
rect 8536 17184 8542 17196
rect 9677 17187 9735 17193
rect 9677 17184 9689 17187
rect 8536 17156 9689 17184
rect 8536 17144 8542 17156
rect 9677 17153 9689 17156
rect 9723 17153 9735 17187
rect 9677 17147 9735 17153
rect 2593 17119 2651 17125
rect 2593 17085 2605 17119
rect 2639 17085 2651 17119
rect 2593 17079 2651 17085
rect 4249 17119 4307 17125
rect 4249 17085 4261 17119
rect 4295 17085 4307 17119
rect 4249 17079 4307 17085
rect 2608 16980 2636 17079
rect 2958 16980 2964 16992
rect 2608 16952 2964 16980
rect 2958 16940 2964 16952
rect 3016 16980 3022 16992
rect 4264 16980 4292 17079
rect 5626 17076 5632 17128
rect 5684 17076 5690 17128
rect 7742 17076 7748 17128
rect 7800 17076 7806 17128
rect 8386 17076 8392 17128
rect 8444 17116 8450 17128
rect 9493 17119 9551 17125
rect 9493 17116 9505 17119
rect 8444 17088 9505 17116
rect 8444 17076 8450 17088
rect 9493 17085 9505 17088
rect 9539 17116 9551 17119
rect 10060 17116 10088 17224
rect 10870 17212 10876 17224
rect 10928 17212 10934 17264
rect 14476 17252 14504 17280
rect 15102 17252 15108 17264
rect 14476 17224 15108 17252
rect 15102 17212 15108 17224
rect 15160 17212 15166 17264
rect 10413 17187 10471 17193
rect 10413 17184 10425 17187
rect 9539 17088 10088 17116
rect 10152 17156 10425 17184
rect 9539 17085 9551 17088
rect 9493 17079 9551 17085
rect 5644 17048 5672 17076
rect 10152 17057 10180 17156
rect 10413 17153 10425 17156
rect 10459 17153 10471 17187
rect 10413 17147 10471 17153
rect 11330 17076 11336 17128
rect 11388 17076 11394 17128
rect 13170 17076 13176 17128
rect 13228 17116 13234 17128
rect 14277 17119 14335 17125
rect 14277 17116 14289 17119
rect 13228 17088 14289 17116
rect 13228 17076 13234 17088
rect 14277 17085 14289 17088
rect 14323 17085 14335 17119
rect 14277 17079 14335 17085
rect 6365 17051 6423 17057
rect 6365 17048 6377 17051
rect 5644 17020 6377 17048
rect 6365 17017 6377 17020
rect 6411 17017 6423 17051
rect 6365 17011 6423 17017
rect 10137 17051 10195 17057
rect 10137 17017 10149 17051
rect 10183 17017 10195 17051
rect 10137 17011 10195 17017
rect 3016 16952 4292 16980
rect 3016 16940 3022 16952
rect 5534 16940 5540 16992
rect 5592 16980 5598 16992
rect 5629 16983 5687 16989
rect 5629 16980 5641 16983
rect 5592 16952 5641 16980
rect 5592 16940 5598 16952
rect 5629 16949 5641 16952
rect 5675 16949 5687 16983
rect 5629 16943 5687 16949
rect 10686 16940 10692 16992
rect 10744 16940 10750 16992
rect 1104 16890 18124 16912
rect 1104 16838 3077 16890
rect 3129 16838 3141 16890
rect 3193 16838 3205 16890
rect 3257 16838 3269 16890
rect 3321 16838 3333 16890
rect 3385 16838 7332 16890
rect 7384 16838 7396 16890
rect 7448 16838 7460 16890
rect 7512 16838 7524 16890
rect 7576 16838 7588 16890
rect 7640 16838 11587 16890
rect 11639 16838 11651 16890
rect 11703 16838 11715 16890
rect 11767 16838 11779 16890
rect 11831 16838 11843 16890
rect 11895 16838 15842 16890
rect 15894 16838 15906 16890
rect 15958 16838 15970 16890
rect 16022 16838 16034 16890
rect 16086 16838 16098 16890
rect 16150 16838 18124 16890
rect 1104 16816 18124 16838
rect 2866 16736 2872 16788
rect 2924 16776 2930 16788
rect 2961 16779 3019 16785
rect 2961 16776 2973 16779
rect 2924 16748 2973 16776
rect 2924 16736 2930 16748
rect 2961 16745 2973 16748
rect 3007 16745 3019 16779
rect 2961 16739 3019 16745
rect 4709 16779 4767 16785
rect 4709 16745 4721 16779
rect 4755 16776 4767 16779
rect 5074 16776 5080 16788
rect 4755 16748 5080 16776
rect 4755 16745 4767 16748
rect 4709 16739 4767 16745
rect 5074 16736 5080 16748
rect 5132 16736 5138 16788
rect 8662 16776 8668 16788
rect 5460 16748 8668 16776
rect 1673 16643 1731 16649
rect 1673 16609 1685 16643
rect 1719 16640 1731 16643
rect 2498 16640 2504 16652
rect 1719 16612 2504 16640
rect 1719 16609 1731 16612
rect 1673 16603 1731 16609
rect 2498 16600 2504 16612
rect 2556 16600 2562 16652
rect 4430 16600 4436 16652
rect 4488 16600 4494 16652
rect 5166 16600 5172 16652
rect 5224 16600 5230 16652
rect 5353 16643 5411 16649
rect 5353 16609 5365 16643
rect 5399 16640 5411 16643
rect 5460 16640 5488 16748
rect 8662 16736 8668 16748
rect 8720 16736 8726 16788
rect 11054 16776 11060 16788
rect 10336 16748 11060 16776
rect 8297 16711 8355 16717
rect 8297 16677 8309 16711
rect 8343 16708 8355 16711
rect 8343 16680 9536 16708
rect 8343 16677 8355 16680
rect 8297 16671 8355 16677
rect 5399 16612 5488 16640
rect 5399 16609 5411 16612
rect 5353 16603 5411 16609
rect 5534 16600 5540 16652
rect 5592 16640 5598 16652
rect 9508 16649 9536 16680
rect 6089 16643 6147 16649
rect 6089 16640 6101 16643
rect 5592 16612 6101 16640
rect 5592 16600 5598 16612
rect 6089 16609 6101 16612
rect 6135 16609 6147 16643
rect 6089 16603 6147 16609
rect 9493 16643 9551 16649
rect 9493 16609 9505 16643
rect 9539 16640 9551 16643
rect 9582 16640 9588 16652
rect 9539 16612 9588 16640
rect 9539 16609 9551 16612
rect 9493 16603 9551 16609
rect 9582 16600 9588 16612
rect 9640 16600 9646 16652
rect 10336 16649 10364 16748
rect 11054 16736 11060 16748
rect 11112 16736 11118 16788
rect 11330 16736 11336 16788
rect 11388 16776 11394 16788
rect 11701 16779 11759 16785
rect 11701 16776 11713 16779
rect 11388 16748 11713 16776
rect 11388 16736 11394 16748
rect 11701 16745 11713 16748
rect 11747 16776 11759 16779
rect 11747 16748 12434 16776
rect 11747 16745 11759 16748
rect 11701 16739 11759 16745
rect 12406 16708 12434 16748
rect 15473 16711 15531 16717
rect 12406 16680 12664 16708
rect 10321 16643 10379 16649
rect 10321 16609 10333 16643
rect 10367 16609 10379 16643
rect 10321 16603 10379 16609
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16640 11943 16643
rect 11974 16640 11980 16652
rect 11931 16612 11980 16640
rect 11931 16609 11943 16612
rect 11885 16603 11943 16609
rect 11974 16600 11980 16612
rect 12032 16600 12038 16652
rect 12526 16600 12532 16652
rect 12584 16600 12590 16652
rect 12636 16640 12664 16680
rect 15473 16677 15485 16711
rect 15519 16677 15531 16711
rect 15473 16671 15531 16677
rect 12894 16640 12900 16652
rect 12952 16649 12958 16652
rect 12952 16643 12980 16649
rect 12636 16612 12900 16640
rect 12894 16600 12900 16612
rect 12968 16609 12980 16643
rect 12952 16603 12980 16609
rect 12952 16600 12958 16603
rect 13078 16600 13084 16652
rect 13136 16600 13142 16652
rect 13725 16643 13783 16649
rect 13725 16609 13737 16643
rect 13771 16640 13783 16643
rect 14458 16640 14464 16652
rect 13771 16612 14464 16640
rect 13771 16609 13783 16612
rect 13725 16603 13783 16609
rect 14458 16600 14464 16612
rect 14516 16600 14522 16652
rect 3145 16575 3203 16581
rect 3145 16541 3157 16575
rect 3191 16572 3203 16575
rect 3191 16544 3832 16572
rect 3191 16541 3203 16544
rect 3145 16535 3203 16541
rect 842 16464 848 16516
rect 900 16504 906 16516
rect 1489 16507 1547 16513
rect 1489 16504 1501 16507
rect 900 16476 1501 16504
rect 900 16464 906 16476
rect 1489 16473 1501 16476
rect 1535 16473 1547 16507
rect 1489 16467 1547 16473
rect 3804 16445 3832 16544
rect 4154 16532 4160 16584
rect 4212 16532 4218 16584
rect 4246 16532 4252 16584
rect 4304 16572 4310 16584
rect 5184 16572 5212 16600
rect 4304 16544 5212 16572
rect 4304 16532 4310 16544
rect 6914 16532 6920 16584
rect 6972 16572 6978 16584
rect 7742 16572 7748 16584
rect 6972 16544 7748 16572
rect 6972 16532 6978 16544
rect 7742 16532 7748 16544
rect 7800 16532 7806 16584
rect 8754 16532 8760 16584
rect 8812 16572 8818 16584
rect 10226 16572 10232 16584
rect 8812 16544 10232 16572
rect 8812 16532 8818 16544
rect 10226 16532 10232 16544
rect 10284 16532 10290 16584
rect 10870 16532 10876 16584
rect 10928 16572 10934 16584
rect 11606 16572 11612 16584
rect 10928 16544 11612 16572
rect 10928 16532 10934 16544
rect 11606 16532 11612 16544
rect 11664 16532 11670 16584
rect 12066 16532 12072 16584
rect 12124 16532 12130 16584
rect 12802 16532 12808 16584
rect 12860 16532 12866 16584
rect 15286 16532 15292 16584
rect 15344 16532 15350 16584
rect 7190 16513 7196 16516
rect 5077 16507 5135 16513
rect 5077 16473 5089 16507
rect 5123 16504 5135 16507
rect 5537 16507 5595 16513
rect 5537 16504 5549 16507
rect 5123 16476 5549 16504
rect 5123 16473 5135 16476
rect 5077 16467 5135 16473
rect 5537 16473 5549 16476
rect 5583 16473 5595 16507
rect 5537 16467 5595 16473
rect 7184 16467 7196 16513
rect 7190 16464 7196 16467
rect 7248 16464 7254 16516
rect 9214 16504 9220 16516
rect 8404 16476 9220 16504
rect 3789 16439 3847 16445
rect 3789 16405 3801 16439
rect 3835 16405 3847 16439
rect 3789 16399 3847 16405
rect 5442 16396 5448 16448
rect 5500 16436 5506 16448
rect 8404 16436 8432 16476
rect 9214 16464 9220 16476
rect 9272 16464 9278 16516
rect 10588 16507 10646 16513
rect 10588 16473 10600 16507
rect 10634 16504 10646 16507
rect 11514 16504 11520 16516
rect 10634 16476 11520 16504
rect 10634 16473 10646 16476
rect 10588 16467 10646 16473
rect 11514 16464 11520 16476
rect 11572 16464 11578 16516
rect 15488 16504 15516 16671
rect 15562 16600 15568 16652
rect 15620 16600 15626 16652
rect 17589 16575 17647 16581
rect 17589 16572 17601 16575
rect 16960 16544 17601 16572
rect 15810 16507 15868 16513
rect 15810 16504 15822 16507
rect 15488 16476 15822 16504
rect 15810 16473 15822 16476
rect 15856 16473 15868 16507
rect 15810 16467 15868 16473
rect 5500 16408 8432 16436
rect 5500 16396 5506 16408
rect 8938 16396 8944 16448
rect 8996 16396 9002 16448
rect 12066 16396 12072 16448
rect 12124 16436 12130 16448
rect 16960 16445 16988 16544
rect 17589 16541 17601 16544
rect 17635 16541 17647 16575
rect 17589 16535 17647 16541
rect 16945 16439 17003 16445
rect 16945 16436 16957 16439
rect 12124 16408 16957 16436
rect 12124 16396 12130 16408
rect 16945 16405 16957 16408
rect 16991 16405 17003 16439
rect 16945 16399 17003 16405
rect 17034 16396 17040 16448
rect 17092 16396 17098 16448
rect 1104 16346 18124 16368
rect 1104 16294 3737 16346
rect 3789 16294 3801 16346
rect 3853 16294 3865 16346
rect 3917 16294 3929 16346
rect 3981 16294 3993 16346
rect 4045 16294 7992 16346
rect 8044 16294 8056 16346
rect 8108 16294 8120 16346
rect 8172 16294 8184 16346
rect 8236 16294 8248 16346
rect 8300 16294 12247 16346
rect 12299 16294 12311 16346
rect 12363 16294 12375 16346
rect 12427 16294 12439 16346
rect 12491 16294 12503 16346
rect 12555 16294 16502 16346
rect 16554 16294 16566 16346
rect 16618 16294 16630 16346
rect 16682 16294 16694 16346
rect 16746 16294 16758 16346
rect 16810 16294 18124 16346
rect 1104 16272 18124 16294
rect 7190 16192 7196 16244
rect 7248 16192 7254 16244
rect 7837 16235 7895 16241
rect 7837 16201 7849 16235
rect 7883 16232 7895 16235
rect 8938 16232 8944 16244
rect 7883 16204 8944 16232
rect 7883 16201 7895 16204
rect 7837 16195 7895 16201
rect 8938 16192 8944 16204
rect 8996 16192 9002 16244
rect 9214 16192 9220 16244
rect 9272 16232 9278 16244
rect 10594 16232 10600 16244
rect 9272 16204 10600 16232
rect 9272 16192 9278 16204
rect 10594 16192 10600 16204
rect 10652 16192 10658 16244
rect 10686 16192 10692 16244
rect 10744 16232 10750 16244
rect 10965 16235 11023 16241
rect 10965 16232 10977 16235
rect 10744 16204 10977 16232
rect 10744 16192 10750 16204
rect 10965 16201 10977 16204
rect 11011 16201 11023 16235
rect 10965 16195 11023 16201
rect 11333 16235 11391 16241
rect 11333 16201 11345 16235
rect 11379 16201 11391 16235
rect 11333 16195 11391 16201
rect 4430 16124 4436 16176
rect 4488 16164 4494 16176
rect 8754 16164 8760 16176
rect 4488 16136 8760 16164
rect 4488 16124 4494 16136
rect 2958 16056 2964 16108
rect 3016 16096 3022 16108
rect 3418 16105 3424 16108
rect 3145 16099 3203 16105
rect 3145 16096 3157 16099
rect 3016 16068 3157 16096
rect 3016 16056 3022 16068
rect 3145 16065 3157 16068
rect 3191 16065 3203 16099
rect 3145 16059 3203 16065
rect 3412 16059 3424 16105
rect 3418 16056 3424 16059
rect 3476 16056 3482 16108
rect 5169 16099 5227 16105
rect 5169 16096 5181 16099
rect 4540 16068 5181 16096
rect 4540 15969 4568 16068
rect 5169 16065 5181 16068
rect 5215 16096 5227 16099
rect 5350 16096 5356 16108
rect 5215 16068 5356 16096
rect 5215 16065 5227 16068
rect 5169 16059 5227 16065
rect 5350 16056 5356 16068
rect 5408 16096 5414 16108
rect 5810 16096 5816 16108
rect 5408 16068 5816 16096
rect 5408 16056 5414 16068
rect 5810 16056 5816 16068
rect 5868 16056 5874 16108
rect 7377 16099 7435 16105
rect 7377 16065 7389 16099
rect 7423 16096 7435 16099
rect 7423 16068 7512 16096
rect 7423 16065 7435 16068
rect 7377 16059 7435 16065
rect 4525 15963 4583 15969
rect 4525 15929 4537 15963
rect 4571 15929 4583 15963
rect 4525 15923 4583 15929
rect 5258 15920 5264 15972
rect 5316 15960 5322 15972
rect 5718 15960 5724 15972
rect 5316 15932 5724 15960
rect 5316 15920 5322 15932
rect 5718 15920 5724 15932
rect 5776 15920 5782 15972
rect 7484 15969 7512 16068
rect 7834 15988 7840 16040
rect 7892 16028 7898 16040
rect 8036 16037 8064 16136
rect 8754 16124 8760 16136
rect 8812 16124 8818 16176
rect 10873 16167 10931 16173
rect 10873 16133 10885 16167
rect 10919 16164 10931 16167
rect 11146 16164 11152 16176
rect 10919 16136 11152 16164
rect 10919 16133 10931 16136
rect 10873 16127 10931 16133
rect 11146 16124 11152 16136
rect 11204 16124 11210 16176
rect 8573 16099 8631 16105
rect 8573 16065 8585 16099
rect 8619 16096 8631 16099
rect 8619 16068 8984 16096
rect 8619 16065 8631 16068
rect 8573 16059 8631 16065
rect 8956 16040 8984 16068
rect 9582 16056 9588 16108
rect 9640 16105 9646 16108
rect 9640 16099 9668 16105
rect 9656 16065 9668 16099
rect 10704 16096 10824 16100
rect 11348 16096 11376 16195
rect 11514 16192 11520 16244
rect 11572 16192 11578 16244
rect 11606 16192 11612 16244
rect 11664 16232 11670 16244
rect 11664 16204 14688 16232
rect 11664 16192 11670 16204
rect 11701 16099 11759 16105
rect 11701 16096 11713 16099
rect 9640 16059 9668 16065
rect 10428 16072 11284 16096
rect 10428 16068 10732 16072
rect 10796 16068 11284 16072
rect 11348 16068 11713 16096
rect 9640 16056 9646 16059
rect 7929 16031 7987 16037
rect 7929 16028 7941 16031
rect 7892 16000 7941 16028
rect 7892 15988 7898 16000
rect 7929 15997 7941 16000
rect 7975 15997 7987 16031
rect 7929 15991 7987 15997
rect 8021 16031 8079 16037
rect 8021 15997 8033 16031
rect 8067 15997 8079 16031
rect 8021 15991 8079 15997
rect 8757 16031 8815 16037
rect 8757 15997 8769 16031
rect 8803 15997 8815 16031
rect 8757 15991 8815 15997
rect 7469 15963 7527 15969
rect 7469 15929 7481 15963
rect 7515 15929 7527 15963
rect 7469 15923 7527 15929
rect 4614 15852 4620 15904
rect 4672 15852 4678 15904
rect 4706 15852 4712 15904
rect 4764 15892 4770 15904
rect 6086 15892 6092 15904
rect 4764 15864 6092 15892
rect 4764 15852 4770 15864
rect 6086 15852 6092 15864
rect 6144 15852 6150 15904
rect 8772 15892 8800 15991
rect 8938 15988 8944 16040
rect 8996 16028 9002 16040
rect 9306 16028 9312 16040
rect 8996 16000 9312 16028
rect 8996 15988 9002 16000
rect 9306 15988 9312 16000
rect 9364 15988 9370 16040
rect 9490 15988 9496 16040
rect 9548 15988 9554 16040
rect 9769 16031 9827 16037
rect 9769 15997 9781 16031
rect 9815 16028 9827 16031
rect 9950 16028 9956 16040
rect 9815 16000 9956 16028
rect 9815 15997 9827 16000
rect 9769 15991 9827 15997
rect 9950 15988 9956 16000
rect 10008 16028 10014 16040
rect 10428 16028 10456 16068
rect 10008 16000 10456 16028
rect 10781 16031 10839 16037
rect 10008 15988 10014 16000
rect 10781 15997 10793 16031
rect 10827 15997 10839 16031
rect 11256 16028 11284 16068
rect 11701 16065 11713 16068
rect 11747 16065 11759 16099
rect 11701 16059 11759 16065
rect 11882 16056 11888 16108
rect 11940 16056 11946 16108
rect 12066 16056 12072 16108
rect 12124 16056 12130 16108
rect 12802 16056 12808 16108
rect 12860 16056 12866 16108
rect 12894 16056 12900 16108
rect 12952 16105 12958 16108
rect 12952 16099 12980 16105
rect 12968 16065 12980 16099
rect 12952 16059 12980 16065
rect 12952 16056 12958 16059
rect 13081 16031 13139 16037
rect 13081 16028 13093 16031
rect 11256 16000 13093 16028
rect 10781 15991 10839 15997
rect 13081 15997 13093 16000
rect 13127 16028 13139 16031
rect 13127 16000 14605 16028
rect 13127 15997 13139 16000
rect 13081 15991 13139 15997
rect 9214 15920 9220 15972
rect 9272 15920 9278 15972
rect 10226 15920 10232 15972
rect 10284 15960 10290 15972
rect 10686 15960 10692 15972
rect 10284 15932 10692 15960
rect 10284 15920 10290 15932
rect 10686 15920 10692 15932
rect 10744 15960 10750 15972
rect 10796 15960 10824 15991
rect 12526 15960 12532 15972
rect 10744 15932 10824 15960
rect 12452 15932 12532 15960
rect 10744 15920 10750 15932
rect 9122 15892 9128 15904
rect 8772 15864 9128 15892
rect 9122 15852 9128 15864
rect 9180 15892 9186 15904
rect 10134 15892 10140 15904
rect 9180 15864 10140 15892
rect 9180 15852 9186 15864
rect 10134 15852 10140 15864
rect 10192 15852 10198 15904
rect 10318 15852 10324 15904
rect 10376 15892 10382 15904
rect 10413 15895 10471 15901
rect 10413 15892 10425 15895
rect 10376 15864 10425 15892
rect 10376 15852 10382 15864
rect 10413 15861 10425 15864
rect 10459 15861 10471 15895
rect 10413 15855 10471 15861
rect 10594 15852 10600 15904
rect 10652 15892 10658 15904
rect 12452 15892 12480 15932
rect 12526 15920 12532 15932
rect 12584 15920 12590 15972
rect 10652 15864 12480 15892
rect 10652 15852 10658 15864
rect 13262 15852 13268 15904
rect 13320 15892 13326 15904
rect 13725 15895 13783 15901
rect 13725 15892 13737 15895
rect 13320 15864 13737 15892
rect 13320 15852 13326 15864
rect 13725 15861 13737 15864
rect 13771 15861 13783 15895
rect 14577 15892 14605 16000
rect 14660 15960 14688 16204
rect 15286 16192 15292 16244
rect 15344 16232 15350 16244
rect 15473 16235 15531 16241
rect 15473 16232 15485 16235
rect 15344 16204 15485 16232
rect 15344 16192 15350 16204
rect 15473 16201 15485 16204
rect 15519 16201 15531 16235
rect 15473 16195 15531 16201
rect 15841 16235 15899 16241
rect 15841 16201 15853 16235
rect 15887 16232 15899 16235
rect 17034 16232 17040 16244
rect 15887 16204 17040 16232
rect 15887 16201 15899 16204
rect 15841 16195 15899 16201
rect 17034 16192 17040 16204
rect 17092 16192 17098 16244
rect 14918 16124 14924 16176
rect 14976 16164 14982 16176
rect 15933 16167 15991 16173
rect 15933 16164 15945 16167
rect 14976 16136 15945 16164
rect 14976 16124 14982 16136
rect 15933 16133 15945 16136
rect 15979 16133 15991 16167
rect 15933 16127 15991 16133
rect 15194 16056 15200 16108
rect 15252 16096 15258 16108
rect 17497 16099 17555 16105
rect 17497 16096 17509 16099
rect 15252 16068 17509 16096
rect 15252 16056 15258 16068
rect 17497 16065 17509 16068
rect 17543 16065 17555 16099
rect 17497 16059 17555 16065
rect 16025 16031 16083 16037
rect 16025 15997 16037 16031
rect 16071 15997 16083 16031
rect 16025 15991 16083 15997
rect 15654 15960 15660 15972
rect 14660 15932 15660 15960
rect 15654 15920 15660 15932
rect 15712 15960 15718 15972
rect 16040 15960 16068 15991
rect 16482 15988 16488 16040
rect 16540 16028 16546 16040
rect 17221 16031 17279 16037
rect 17221 16028 17233 16031
rect 16540 16000 17233 16028
rect 16540 15988 16546 16000
rect 17221 15997 17233 16000
rect 17267 15997 17279 16031
rect 17221 15991 17279 15997
rect 15712 15932 16068 15960
rect 15712 15920 15718 15932
rect 14734 15892 14740 15904
rect 14577 15864 14740 15892
rect 13725 15855 13783 15861
rect 14734 15852 14740 15864
rect 14792 15852 14798 15904
rect 15746 15852 15752 15904
rect 15804 15892 15810 15904
rect 16669 15895 16727 15901
rect 16669 15892 16681 15895
rect 15804 15864 16681 15892
rect 15804 15852 15810 15864
rect 16669 15861 16681 15864
rect 16715 15861 16727 15895
rect 16669 15855 16727 15861
rect 17678 15852 17684 15904
rect 17736 15852 17742 15904
rect 1104 15802 18124 15824
rect 1104 15750 3077 15802
rect 3129 15750 3141 15802
rect 3193 15750 3205 15802
rect 3257 15750 3269 15802
rect 3321 15750 3333 15802
rect 3385 15750 7332 15802
rect 7384 15750 7396 15802
rect 7448 15750 7460 15802
rect 7512 15750 7524 15802
rect 7576 15750 7588 15802
rect 7640 15750 11587 15802
rect 11639 15750 11651 15802
rect 11703 15750 11715 15802
rect 11767 15750 11779 15802
rect 11831 15750 11843 15802
rect 11895 15750 15842 15802
rect 15894 15750 15906 15802
rect 15958 15750 15970 15802
rect 16022 15750 16034 15802
rect 16086 15750 16098 15802
rect 16150 15750 18124 15802
rect 1104 15728 18124 15750
rect 3418 15648 3424 15700
rect 3476 15648 3482 15700
rect 4706 15688 4712 15700
rect 3712 15660 4712 15688
rect 3712 15620 3740 15660
rect 4706 15648 4712 15660
rect 4764 15648 4770 15700
rect 5534 15688 5540 15700
rect 4816 15660 5540 15688
rect 1688 15592 3740 15620
rect 3789 15623 3847 15629
rect 1688 15493 1716 15592
rect 3789 15589 3801 15623
rect 3835 15589 3847 15623
rect 3789 15583 3847 15589
rect 2498 15512 2504 15564
rect 2556 15552 2562 15564
rect 2556 15524 2774 15552
rect 2556 15512 2562 15524
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15453 1731 15487
rect 1673 15447 1731 15453
rect 2746 15416 2774 15524
rect 3605 15487 3663 15493
rect 3605 15453 3617 15487
rect 3651 15484 3663 15487
rect 3804 15484 3832 15583
rect 4246 15512 4252 15564
rect 4304 15512 4310 15564
rect 4430 15512 4436 15564
rect 4488 15512 4494 15564
rect 3651 15456 3832 15484
rect 4157 15487 4215 15493
rect 3651 15453 3663 15456
rect 3605 15447 3663 15453
rect 4157 15453 4169 15487
rect 4203 15484 4215 15487
rect 4614 15484 4620 15496
rect 4203 15456 4620 15484
rect 4203 15453 4215 15456
rect 4157 15447 4215 15453
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 4706 15444 4712 15496
rect 4764 15484 4770 15496
rect 4816 15493 4844 15660
rect 5534 15648 5540 15660
rect 5592 15648 5598 15700
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 9858 15688 9864 15700
rect 9548 15660 9864 15688
rect 9548 15648 9554 15660
rect 9858 15648 9864 15660
rect 9916 15648 9922 15700
rect 5442 15552 5448 15564
rect 5184 15524 5448 15552
rect 5184 15496 5212 15524
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 5810 15512 5816 15564
rect 5868 15561 5874 15564
rect 5868 15555 5896 15561
rect 5884 15521 5896 15555
rect 5868 15515 5896 15521
rect 5997 15555 6055 15561
rect 5997 15521 6009 15555
rect 6043 15552 6055 15555
rect 7098 15552 7104 15564
rect 6043 15524 7104 15552
rect 6043 15521 6055 15524
rect 5997 15515 6055 15521
rect 5868 15512 5874 15515
rect 7098 15512 7104 15524
rect 7156 15512 7162 15564
rect 8938 15512 8944 15564
rect 8996 15512 9002 15564
rect 9122 15512 9128 15564
rect 9180 15512 9186 15564
rect 9585 15555 9643 15561
rect 9585 15552 9597 15555
rect 9232 15524 9597 15552
rect 4801 15487 4859 15493
rect 4801 15484 4813 15487
rect 4764 15456 4813 15484
rect 4764 15444 4770 15456
rect 4801 15453 4813 15456
rect 4847 15453 4859 15487
rect 4801 15447 4859 15453
rect 4890 15444 4896 15496
rect 4948 15484 4954 15496
rect 4985 15487 5043 15493
rect 4985 15484 4997 15487
rect 4948 15456 4997 15484
rect 4948 15444 4954 15456
rect 4985 15453 4997 15456
rect 5031 15453 5043 15487
rect 4985 15447 5043 15453
rect 4246 15416 4252 15428
rect 2746 15388 4252 15416
rect 4246 15376 4252 15388
rect 4304 15376 4310 15428
rect 1486 15308 1492 15360
rect 1544 15308 1550 15360
rect 5000 15348 5028 15447
rect 5166 15444 5172 15496
rect 5224 15444 5230 15496
rect 5718 15444 5724 15496
rect 5776 15444 5782 15496
rect 7469 15487 7527 15493
rect 7469 15453 7481 15487
rect 7515 15484 7527 15487
rect 7650 15484 7656 15496
rect 7515 15456 7656 15484
rect 7515 15453 7527 15456
rect 7469 15447 7527 15453
rect 7650 15444 7656 15456
rect 7708 15444 7714 15496
rect 9232 15484 9260 15524
rect 9585 15521 9597 15524
rect 9631 15521 9643 15555
rect 9585 15515 9643 15521
rect 9674 15512 9680 15564
rect 9732 15552 9738 15564
rect 9978 15555 10036 15561
rect 9978 15552 9990 15555
rect 9732 15524 9990 15552
rect 9732 15512 9738 15524
rect 9978 15521 9990 15524
rect 10024 15521 10036 15555
rect 9978 15515 10036 15521
rect 10137 15555 10195 15561
rect 10137 15521 10149 15555
rect 10183 15552 10195 15555
rect 10183 15524 12434 15552
rect 10183 15521 10195 15524
rect 10137 15515 10195 15521
rect 9140 15456 9260 15484
rect 9140 15416 9168 15456
rect 9858 15444 9864 15496
rect 9916 15444 9922 15496
rect 12406 15484 12434 15524
rect 12526 15512 12532 15564
rect 12584 15552 12590 15564
rect 15289 15555 15347 15561
rect 15289 15552 15301 15555
rect 12584 15524 15301 15552
rect 12584 15512 12590 15524
rect 15289 15521 15301 15524
rect 15335 15521 15347 15555
rect 15289 15515 15347 15521
rect 15562 15512 15568 15564
rect 15620 15552 15626 15564
rect 16025 15555 16083 15561
rect 16025 15552 16037 15555
rect 15620 15524 16037 15552
rect 15620 15512 15626 15524
rect 16025 15521 16037 15524
rect 16071 15521 16083 15555
rect 16025 15515 16083 15521
rect 12710 15484 12716 15496
rect 12406 15456 12716 15484
rect 12710 15444 12716 15456
rect 12768 15484 12774 15496
rect 13078 15484 13084 15496
rect 12768 15456 13084 15484
rect 12768 15444 12774 15456
rect 13078 15444 13084 15456
rect 13136 15444 13142 15496
rect 13173 15487 13231 15493
rect 13173 15453 13185 15487
rect 13219 15484 13231 15487
rect 13906 15484 13912 15496
rect 13219 15456 13912 15484
rect 13219 15453 13231 15456
rect 13173 15447 13231 15453
rect 13906 15444 13912 15456
rect 13964 15444 13970 15496
rect 14734 15444 14740 15496
rect 14792 15444 14798 15496
rect 14826 15444 14832 15496
rect 14884 15493 14890 15496
rect 14884 15487 14933 15493
rect 14884 15453 14887 15487
rect 14921 15453 14933 15487
rect 14884 15447 14933 15453
rect 14884 15444 14890 15447
rect 15010 15444 15016 15496
rect 15068 15444 15074 15496
rect 15749 15487 15807 15493
rect 15749 15453 15761 15487
rect 15795 15484 15807 15487
rect 15838 15484 15844 15496
rect 15795 15456 15844 15484
rect 15795 15453 15807 15456
rect 15749 15447 15807 15453
rect 15838 15444 15844 15456
rect 15896 15444 15902 15496
rect 15933 15487 15991 15493
rect 15933 15453 15945 15487
rect 15979 15484 15991 15487
rect 16114 15484 16120 15496
rect 15979 15456 16120 15484
rect 15979 15453 15991 15456
rect 15933 15447 15991 15453
rect 16114 15444 16120 15456
rect 16172 15444 16178 15496
rect 17494 15444 17500 15496
rect 17552 15444 17558 15496
rect 12802 15416 12808 15428
rect 6564 15388 9168 15416
rect 5626 15348 5632 15360
rect 5000 15320 5632 15348
rect 5626 15308 5632 15320
rect 5684 15308 5690 15360
rect 5718 15308 5724 15360
rect 5776 15348 5782 15360
rect 6564 15348 6592 15388
rect 5776 15320 6592 15348
rect 5776 15308 5782 15320
rect 6638 15308 6644 15360
rect 6696 15308 6702 15360
rect 7282 15308 7288 15360
rect 7340 15308 7346 15360
rect 9140 15348 9168 15388
rect 10612 15388 12808 15416
rect 10612 15348 10640 15388
rect 12802 15376 12808 15388
rect 12860 15416 12866 15428
rect 13722 15416 13728 15428
rect 12860 15388 13728 15416
rect 12860 15376 12866 15388
rect 13722 15376 13728 15388
rect 13780 15376 13786 15428
rect 16298 15425 16304 15428
rect 16292 15379 16304 15425
rect 16298 15376 16304 15379
rect 16356 15376 16362 15428
rect 9140 15320 10640 15348
rect 10778 15308 10784 15360
rect 10836 15308 10842 15360
rect 12529 15351 12587 15357
rect 12529 15317 12541 15351
rect 12575 15348 12587 15351
rect 12618 15348 12624 15360
rect 12575 15320 12624 15348
rect 12575 15317 12587 15320
rect 12529 15311 12587 15317
rect 12618 15308 12624 15320
rect 12676 15308 12682 15360
rect 14093 15351 14151 15357
rect 14093 15317 14105 15351
rect 14139 15348 14151 15351
rect 14274 15348 14280 15360
rect 14139 15320 14280 15348
rect 14139 15317 14151 15320
rect 14093 15311 14151 15317
rect 14274 15308 14280 15320
rect 14332 15308 14338 15360
rect 15838 15308 15844 15360
rect 15896 15348 15902 15360
rect 16482 15348 16488 15360
rect 15896 15320 16488 15348
rect 15896 15308 15902 15320
rect 16482 15308 16488 15320
rect 16540 15348 16546 15360
rect 17405 15351 17463 15357
rect 17405 15348 17417 15351
rect 16540 15320 17417 15348
rect 16540 15308 16546 15320
rect 17405 15317 17417 15320
rect 17451 15317 17463 15351
rect 17405 15311 17463 15317
rect 17678 15308 17684 15360
rect 17736 15308 17742 15360
rect 1104 15258 18124 15280
rect 1104 15206 3737 15258
rect 3789 15206 3801 15258
rect 3853 15206 3865 15258
rect 3917 15206 3929 15258
rect 3981 15206 3993 15258
rect 4045 15206 7992 15258
rect 8044 15206 8056 15258
rect 8108 15206 8120 15258
rect 8172 15206 8184 15258
rect 8236 15206 8248 15258
rect 8300 15206 12247 15258
rect 12299 15206 12311 15258
rect 12363 15206 12375 15258
rect 12427 15206 12439 15258
rect 12491 15206 12503 15258
rect 12555 15206 16502 15258
rect 16554 15206 16566 15258
rect 16618 15206 16630 15258
rect 16682 15206 16694 15258
rect 16746 15206 16758 15258
rect 16810 15206 18124 15258
rect 1104 15184 18124 15206
rect 9766 15104 9772 15156
rect 9824 15144 9830 15156
rect 9953 15147 10011 15153
rect 9953 15144 9965 15147
rect 9824 15116 9965 15144
rect 9824 15104 9830 15116
rect 9953 15113 9965 15116
rect 9999 15113 10011 15147
rect 9953 15107 10011 15113
rect 10502 15104 10508 15156
rect 10560 15104 10566 15156
rect 11333 15147 11391 15153
rect 11333 15113 11345 15147
rect 11379 15113 11391 15147
rect 11333 15107 11391 15113
rect 12897 15147 12955 15153
rect 12897 15113 12909 15147
rect 12943 15144 12955 15147
rect 13906 15144 13912 15156
rect 12943 15116 13912 15144
rect 12943 15113 12955 15116
rect 12897 15107 12955 15113
rect 7184 15079 7242 15085
rect 7184 15045 7196 15079
rect 7230 15076 7242 15079
rect 7282 15076 7288 15088
rect 7230 15048 7288 15076
rect 7230 15045 7242 15048
rect 7184 15039 7242 15045
rect 7282 15036 7288 15048
rect 7340 15036 7346 15088
rect 8662 15036 8668 15088
rect 8720 15076 8726 15088
rect 11348 15076 11376 15107
rect 13906 15104 13912 15116
rect 13964 15144 13970 15156
rect 14826 15144 14832 15156
rect 13964 15116 14832 15144
rect 13964 15104 13970 15116
rect 14826 15104 14832 15116
rect 14884 15104 14890 15156
rect 15746 15104 15752 15156
rect 15804 15144 15810 15156
rect 15841 15147 15899 15153
rect 15841 15144 15853 15147
rect 15804 15116 15853 15144
rect 15804 15104 15810 15116
rect 15841 15113 15853 15116
rect 15887 15113 15899 15147
rect 15841 15107 15899 15113
rect 16209 15147 16267 15153
rect 16209 15113 16221 15147
rect 16255 15113 16267 15147
rect 16209 15107 16267 15113
rect 11762 15079 11820 15085
rect 11762 15076 11774 15079
rect 8720 15048 11008 15076
rect 11348 15048 11774 15076
rect 8720 15036 8726 15048
rect 10980 15020 11008 15048
rect 11762 15045 11774 15048
rect 11808 15045 11820 15079
rect 11762 15039 11820 15045
rect 1762 15017 1768 15020
rect 1756 14971 1768 15017
rect 1762 14968 1768 14971
rect 1820 14968 1826 15020
rect 4341 15011 4399 15017
rect 4341 14977 4353 15011
rect 4387 15008 4399 15011
rect 4706 15008 4712 15020
rect 4387 14980 4712 15008
rect 4387 14977 4399 14980
rect 4341 14971 4399 14977
rect 4706 14968 4712 14980
rect 4764 14968 4770 15020
rect 5258 14968 5264 15020
rect 5316 14968 5322 15020
rect 5350 14968 5356 15020
rect 5408 15017 5414 15020
rect 5408 15011 5436 15017
rect 5424 14977 5436 15011
rect 5408 14971 5436 14977
rect 5408 14968 5414 14971
rect 6546 14968 6552 15020
rect 6604 14968 6610 15020
rect 6638 14968 6644 15020
rect 6696 15008 6702 15020
rect 6733 15011 6791 15017
rect 6733 15008 6745 15011
rect 6696 14980 6745 15008
rect 6696 14968 6702 14980
rect 6733 14977 6745 14980
rect 6779 14977 6791 15011
rect 6733 14971 6791 14977
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 8478 15008 8484 15020
rect 6871 14980 8484 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 8478 14968 8484 14980
rect 8536 15008 8542 15020
rect 8536 14980 9260 15008
rect 8536 14968 8542 14980
rect 1394 14900 1400 14952
rect 1452 14940 1458 14952
rect 1489 14943 1547 14949
rect 1489 14940 1501 14943
rect 1452 14912 1501 14940
rect 1452 14900 1458 14912
rect 1489 14909 1501 14912
rect 1535 14909 1547 14943
rect 1489 14903 1547 14909
rect 3513 14943 3571 14949
rect 3513 14909 3525 14943
rect 3559 14909 3571 14943
rect 3513 14903 3571 14909
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14940 4583 14943
rect 4890 14940 4896 14952
rect 4571 14912 4896 14940
rect 4571 14909 4583 14912
rect 4525 14903 4583 14909
rect 2774 14832 2780 14884
rect 2832 14872 2838 14884
rect 2961 14875 3019 14881
rect 2961 14872 2973 14875
rect 2832 14844 2973 14872
rect 2832 14832 2838 14844
rect 2961 14841 2973 14844
rect 3007 14841 3019 14875
rect 2961 14835 3019 14841
rect 3528 14816 3556 14903
rect 4890 14900 4896 14912
rect 4948 14900 4954 14952
rect 5537 14943 5595 14949
rect 5537 14909 5549 14943
rect 5583 14940 5595 14943
rect 5718 14940 5724 14952
rect 5583 14912 5724 14940
rect 5583 14909 5595 14912
rect 5537 14903 5595 14909
rect 5718 14900 5724 14912
rect 5776 14900 5782 14952
rect 6914 14900 6920 14952
rect 6972 14900 6978 14952
rect 8941 14943 8999 14949
rect 8941 14909 8953 14943
rect 8987 14909 8999 14943
rect 9232 14940 9260 14980
rect 9306 14968 9312 15020
rect 9364 14968 9370 15020
rect 10137 15011 10195 15017
rect 10137 14977 10149 15011
rect 10183 15008 10195 15011
rect 10226 15008 10232 15020
rect 10183 14980 10232 15008
rect 10183 14977 10195 14980
rect 10137 14971 10195 14977
rect 10226 14968 10232 14980
rect 10284 14968 10290 15020
rect 10318 14968 10324 15020
rect 10376 14968 10382 15020
rect 10502 14968 10508 15020
rect 10560 15008 10566 15020
rect 10689 15011 10747 15017
rect 10689 15008 10701 15011
rect 10560 14980 10701 15008
rect 10560 14968 10566 14980
rect 10689 14977 10701 14980
rect 10735 14977 10747 15011
rect 10689 14971 10747 14977
rect 10778 14968 10784 15020
rect 10836 15008 10842 15020
rect 10873 15011 10931 15017
rect 10873 15008 10885 15011
rect 10836 14980 10885 15008
rect 10836 14968 10842 14980
rect 10873 14977 10885 14980
rect 10919 14977 10931 15011
rect 10873 14971 10931 14977
rect 10962 14968 10968 15020
rect 11020 14968 11026 15020
rect 11146 14968 11152 15020
rect 11204 14968 11210 15020
rect 13906 15017 13912 15020
rect 13884 15011 13912 15017
rect 13884 14977 13896 15011
rect 13884 14971 13912 14977
rect 13906 14968 13912 14971
rect 13964 14968 13970 15020
rect 15010 15008 15016 15020
rect 14660 14980 15016 15008
rect 10413 14943 10471 14949
rect 10413 14940 10425 14943
rect 9232 14912 10425 14940
rect 8941 14903 8999 14909
rect 10413 14909 10425 14912
rect 10459 14909 10471 14943
rect 10413 14903 10471 14909
rect 4985 14875 5043 14881
rect 4985 14841 4997 14875
rect 5031 14841 5043 14875
rect 4985 14835 5043 14841
rect 8297 14875 8355 14881
rect 8297 14841 8309 14875
rect 8343 14872 8355 14875
rect 8956 14872 8984 14903
rect 10042 14872 10048 14884
rect 8343 14844 10048 14872
rect 8343 14841 8355 14844
rect 8297 14835 8355 14841
rect 2869 14807 2927 14813
rect 2869 14773 2881 14807
rect 2915 14804 2927 14807
rect 3510 14804 3516 14816
rect 2915 14776 3516 14804
rect 2915 14773 2927 14776
rect 2869 14767 2927 14773
rect 3510 14764 3516 14776
rect 3568 14764 3574 14816
rect 5000 14804 5028 14835
rect 10042 14832 10048 14844
rect 10100 14832 10106 14884
rect 5442 14804 5448 14816
rect 5000 14776 5448 14804
rect 5442 14764 5448 14776
rect 5500 14764 5506 14816
rect 6178 14764 6184 14816
rect 6236 14764 6242 14816
rect 6362 14764 6368 14816
rect 6420 14764 6426 14816
rect 8386 14764 8392 14816
rect 8444 14764 8450 14816
rect 9125 14807 9183 14813
rect 9125 14773 9137 14807
rect 9171 14804 9183 14807
rect 9214 14804 9220 14816
rect 9171 14776 9220 14804
rect 9171 14773 9183 14776
rect 9125 14767 9183 14773
rect 9214 14764 9220 14776
rect 9272 14764 9278 14816
rect 10428 14804 10456 14903
rect 11054 14900 11060 14952
rect 11112 14940 11118 14952
rect 11517 14943 11575 14949
rect 11517 14940 11529 14943
rect 11112 14912 11529 14940
rect 11112 14900 11118 14912
rect 11517 14909 11529 14912
rect 11563 14909 11575 14943
rect 11517 14903 11575 14909
rect 12710 14900 12716 14952
rect 12768 14940 12774 14952
rect 13725 14943 13783 14949
rect 13725 14940 13737 14943
rect 12768 14912 13737 14940
rect 12768 14900 12774 14912
rect 13725 14909 13737 14912
rect 13771 14909 13783 14943
rect 13725 14903 13783 14909
rect 14001 14943 14059 14949
rect 14001 14909 14013 14943
rect 14047 14940 14059 14943
rect 14660 14940 14688 14980
rect 15010 14968 15016 14980
rect 15068 14968 15074 15020
rect 16114 15008 16120 15020
rect 15396 14980 16120 15008
rect 14047 14912 14688 14940
rect 14737 14943 14795 14949
rect 14047 14909 14059 14912
rect 14001 14903 14059 14909
rect 14737 14909 14749 14943
rect 14783 14909 14795 14943
rect 14737 14903 14795 14909
rect 14921 14943 14979 14949
rect 14921 14909 14933 14943
rect 14967 14940 14979 14943
rect 15396 14940 15424 14980
rect 16114 14968 16120 14980
rect 16172 14968 16178 15020
rect 16224 15008 16252 15107
rect 16298 15104 16304 15156
rect 16356 15104 16362 15156
rect 16485 15011 16543 15017
rect 16485 15008 16497 15011
rect 16224 14980 16497 15008
rect 16485 14977 16497 14980
rect 16531 14977 16543 15011
rect 16485 14971 16543 14977
rect 17770 14968 17776 15020
rect 17828 14968 17834 15020
rect 14967 14912 15424 14940
rect 14967 14909 14979 14912
rect 14921 14903 14979 14909
rect 14277 14875 14335 14881
rect 14277 14841 14289 14875
rect 14323 14872 14335 14875
rect 14366 14872 14372 14884
rect 14323 14844 14372 14872
rect 14323 14841 14335 14844
rect 14277 14835 14335 14841
rect 14366 14832 14372 14844
rect 14424 14832 14430 14884
rect 14752 14872 14780 14903
rect 15654 14900 15660 14952
rect 15712 14900 15718 14952
rect 15749 14943 15807 14949
rect 15749 14909 15761 14943
rect 15795 14940 15807 14943
rect 15795 14912 15976 14940
rect 15795 14909 15807 14912
rect 15749 14903 15807 14909
rect 15838 14872 15844 14884
rect 14752 14844 15844 14872
rect 15838 14832 15844 14844
rect 15896 14832 15902 14884
rect 12158 14804 12164 14816
rect 10428 14776 12164 14804
rect 12158 14764 12164 14776
rect 12216 14764 12222 14816
rect 13081 14807 13139 14813
rect 13081 14773 13093 14807
rect 13127 14804 13139 14807
rect 14734 14804 14740 14816
rect 13127 14776 14740 14804
rect 13127 14773 13139 14776
rect 13081 14767 13139 14773
rect 14734 14764 14740 14776
rect 14792 14764 14798 14816
rect 15102 14764 15108 14816
rect 15160 14804 15166 14816
rect 15654 14804 15660 14816
rect 15160 14776 15660 14804
rect 15160 14764 15166 14776
rect 15654 14764 15660 14776
rect 15712 14804 15718 14816
rect 15948 14804 15976 14912
rect 16390 14900 16396 14952
rect 16448 14940 16454 14952
rect 17405 14943 17463 14949
rect 17405 14940 17417 14943
rect 16448 14912 17417 14940
rect 16448 14900 16454 14912
rect 17405 14909 17417 14912
rect 17451 14909 17463 14943
rect 17405 14903 17463 14909
rect 15712 14776 15976 14804
rect 15712 14764 15718 14776
rect 16850 14764 16856 14816
rect 16908 14764 16914 14816
rect 17586 14764 17592 14816
rect 17644 14764 17650 14816
rect 1104 14714 18124 14736
rect 1104 14662 3077 14714
rect 3129 14662 3141 14714
rect 3193 14662 3205 14714
rect 3257 14662 3269 14714
rect 3321 14662 3333 14714
rect 3385 14662 7332 14714
rect 7384 14662 7396 14714
rect 7448 14662 7460 14714
rect 7512 14662 7524 14714
rect 7576 14662 7588 14714
rect 7640 14662 11587 14714
rect 11639 14662 11651 14714
rect 11703 14662 11715 14714
rect 11767 14662 11779 14714
rect 11831 14662 11843 14714
rect 11895 14662 15842 14714
rect 15894 14662 15906 14714
rect 15958 14662 15970 14714
rect 16022 14662 16034 14714
rect 16086 14662 16098 14714
rect 16150 14662 18124 14714
rect 1104 14640 18124 14662
rect 1762 14560 1768 14612
rect 1820 14600 1826 14612
rect 1949 14603 2007 14609
rect 1949 14600 1961 14603
rect 1820 14572 1961 14600
rect 1820 14560 1826 14572
rect 1949 14569 1961 14572
rect 1995 14569 2007 14603
rect 1949 14563 2007 14569
rect 6086 14560 6092 14612
rect 6144 14560 6150 14612
rect 6178 14560 6184 14612
rect 6236 14600 6242 14612
rect 6457 14603 6515 14609
rect 6457 14600 6469 14603
rect 6236 14572 6469 14600
rect 6236 14560 6242 14572
rect 6457 14569 6469 14572
rect 6503 14569 6515 14603
rect 6457 14563 6515 14569
rect 10134 14560 10140 14612
rect 10192 14600 10198 14612
rect 10321 14603 10379 14609
rect 10321 14600 10333 14603
rect 10192 14572 10333 14600
rect 10192 14560 10198 14572
rect 10321 14569 10333 14572
rect 10367 14600 10379 14603
rect 10367 14569 10389 14600
rect 10321 14563 10389 14569
rect 842 14492 848 14544
rect 900 14532 906 14544
rect 1489 14535 1547 14541
rect 1489 14532 1501 14535
rect 900 14504 1501 14532
rect 900 14492 906 14504
rect 1489 14501 1501 14504
rect 1535 14501 1547 14535
rect 6362 14532 6368 14544
rect 1489 14495 1547 14501
rect 1964 14504 6368 14532
rect 1673 14399 1731 14405
rect 1673 14365 1685 14399
rect 1719 14396 1731 14399
rect 1964 14396 1992 14504
rect 6362 14492 6368 14504
rect 6420 14492 6426 14544
rect 10361 14532 10389 14563
rect 10962 14560 10968 14612
rect 11020 14600 11026 14612
rect 11020 14572 12434 14600
rect 11020 14560 11026 14572
rect 10361 14504 11008 14532
rect 2314 14424 2320 14476
rect 2372 14464 2378 14476
rect 2869 14467 2927 14473
rect 2869 14464 2881 14467
rect 2372 14436 2881 14464
rect 2372 14424 2378 14436
rect 2869 14433 2881 14436
rect 2915 14433 2927 14467
rect 2869 14427 2927 14433
rect 6549 14467 6607 14473
rect 6549 14433 6561 14467
rect 6595 14464 6607 14467
rect 8662 14464 8668 14476
rect 6595 14436 8668 14464
rect 6595 14433 6607 14436
rect 6549 14427 6607 14433
rect 8662 14424 8668 14436
rect 8720 14424 8726 14476
rect 10980 14473 11008 14504
rect 10965 14467 11023 14473
rect 10965 14433 10977 14467
rect 11011 14433 11023 14467
rect 10965 14427 11023 14433
rect 11054 14424 11060 14476
rect 11112 14464 11118 14476
rect 11330 14464 11336 14476
rect 11112 14436 11336 14464
rect 11112 14424 11118 14436
rect 11330 14424 11336 14436
rect 11388 14464 11394 14476
rect 11885 14467 11943 14473
rect 11885 14464 11897 14467
rect 11388 14436 11897 14464
rect 11388 14424 11394 14436
rect 1719 14368 1992 14396
rect 2133 14399 2191 14405
rect 1719 14365 1731 14368
rect 1673 14359 1731 14365
rect 2133 14365 2145 14399
rect 2179 14396 2191 14399
rect 2685 14399 2743 14405
rect 2179 14368 2360 14396
rect 2179 14365 2191 14368
rect 2133 14359 2191 14365
rect 2332 14269 2360 14368
rect 2685 14365 2697 14399
rect 2731 14396 2743 14399
rect 2774 14396 2780 14408
rect 2731 14368 2780 14396
rect 2731 14365 2743 14368
rect 2685 14359 2743 14365
rect 2774 14356 2780 14368
rect 2832 14356 2838 14408
rect 6270 14356 6276 14408
rect 6328 14356 6334 14408
rect 9214 14405 9220 14408
rect 8941 14399 8999 14405
rect 8941 14396 8953 14399
rect 7024 14368 8953 14396
rect 6914 14288 6920 14340
rect 6972 14328 6978 14340
rect 7024 14337 7052 14368
rect 8941 14365 8953 14368
rect 8987 14365 8999 14399
rect 9208 14396 9220 14405
rect 9175 14368 9220 14396
rect 8941 14359 8999 14365
rect 9208 14359 9220 14368
rect 9214 14356 9220 14359
rect 9272 14356 9278 14408
rect 11624 14405 11652 14436
rect 11885 14433 11897 14436
rect 11931 14433 11943 14467
rect 12406 14464 12434 14572
rect 14090 14560 14096 14612
rect 14148 14560 14154 14612
rect 14458 14560 14464 14612
rect 14516 14560 14522 14612
rect 14734 14560 14740 14612
rect 14792 14560 14798 14612
rect 15105 14603 15163 14609
rect 15105 14569 15117 14603
rect 15151 14600 15163 14603
rect 15194 14600 15200 14612
rect 15151 14572 15200 14600
rect 15151 14569 15163 14572
rect 15105 14563 15163 14569
rect 15194 14560 15200 14572
rect 15252 14560 15258 14612
rect 16301 14603 16359 14609
rect 16301 14569 16313 14603
rect 16347 14600 16359 14603
rect 17770 14600 17776 14612
rect 16347 14572 17776 14600
rect 16347 14569 16359 14572
rect 16301 14563 16359 14569
rect 17770 14560 17776 14572
rect 17828 14560 17834 14612
rect 16390 14492 16396 14544
rect 16448 14492 16454 14544
rect 14553 14467 14611 14473
rect 14553 14464 14565 14467
rect 12406 14436 14565 14464
rect 11885 14427 11943 14433
rect 14553 14433 14565 14436
rect 14599 14464 14611 14467
rect 14645 14467 14703 14473
rect 14645 14464 14657 14467
rect 14599 14436 14657 14464
rect 14599 14433 14611 14436
rect 14553 14427 14611 14433
rect 14645 14433 14657 14436
rect 14691 14433 14703 14467
rect 14645 14427 14703 14433
rect 15746 14424 15752 14476
rect 15804 14424 15810 14476
rect 11609 14399 11667 14405
rect 11609 14365 11621 14399
rect 11655 14396 11667 14399
rect 11655 14368 11689 14396
rect 11655 14365 11667 14368
rect 11609 14359 11667 14365
rect 13446 14356 13452 14408
rect 13504 14396 13510 14408
rect 14277 14399 14335 14405
rect 14277 14396 14289 14399
rect 13504 14368 14289 14396
rect 13504 14356 13510 14368
rect 14277 14365 14289 14368
rect 14323 14365 14335 14399
rect 14277 14359 14335 14365
rect 14366 14356 14372 14408
rect 14424 14396 14430 14408
rect 14921 14399 14979 14405
rect 14921 14396 14933 14399
rect 14424 14368 14933 14396
rect 14424 14356 14430 14368
rect 14921 14365 14933 14368
rect 14967 14365 14979 14399
rect 14921 14359 14979 14365
rect 17506 14399 17564 14405
rect 17506 14365 17518 14399
rect 17552 14365 17564 14399
rect 17506 14359 17564 14365
rect 17773 14399 17831 14405
rect 17773 14365 17785 14399
rect 17819 14365 17831 14399
rect 17773 14359 17831 14365
rect 7009 14331 7067 14337
rect 7009 14328 7021 14331
rect 6972 14300 7021 14328
rect 6972 14288 6978 14300
rect 7009 14297 7021 14300
rect 7055 14297 7067 14331
rect 7009 14291 7067 14297
rect 8754 14288 8760 14340
rect 8812 14288 8818 14340
rect 13633 14331 13691 14337
rect 13633 14297 13645 14331
rect 13679 14328 13691 14331
rect 13722 14328 13728 14340
rect 13679 14300 13728 14328
rect 13679 14297 13691 14300
rect 13633 14291 13691 14297
rect 13722 14288 13728 14300
rect 13780 14288 13786 14340
rect 15654 14288 15660 14340
rect 15712 14328 15718 14340
rect 15841 14331 15899 14337
rect 15841 14328 15853 14331
rect 15712 14300 15853 14328
rect 15712 14288 15718 14300
rect 15841 14297 15853 14300
rect 15887 14297 15899 14331
rect 15841 14291 15899 14297
rect 15933 14331 15991 14337
rect 15933 14297 15945 14331
rect 15979 14328 15991 14331
rect 16850 14328 16856 14340
rect 15979 14300 16856 14328
rect 15979 14297 15991 14300
rect 15933 14291 15991 14297
rect 16850 14288 16856 14300
rect 16908 14288 16914 14340
rect 17512 14328 17540 14359
rect 17586 14328 17592 14340
rect 17512 14300 17592 14328
rect 17586 14288 17592 14300
rect 17644 14288 17650 14340
rect 2317 14263 2375 14269
rect 2317 14229 2329 14263
rect 2363 14229 2375 14263
rect 2317 14223 2375 14229
rect 2498 14220 2504 14272
rect 2556 14260 2562 14272
rect 2777 14263 2835 14269
rect 2777 14260 2789 14263
rect 2556 14232 2789 14260
rect 2556 14220 2562 14232
rect 2777 14229 2789 14232
rect 2823 14229 2835 14263
rect 2777 14223 2835 14229
rect 8938 14220 8944 14272
rect 8996 14260 9002 14272
rect 10413 14263 10471 14269
rect 10413 14260 10425 14263
rect 8996 14232 10425 14260
rect 8996 14220 9002 14232
rect 10413 14229 10425 14232
rect 10459 14229 10471 14263
rect 10413 14223 10471 14229
rect 12066 14220 12072 14272
rect 12124 14260 12130 14272
rect 15470 14260 15476 14272
rect 12124 14232 15476 14260
rect 12124 14220 12130 14232
rect 15470 14220 15476 14232
rect 15528 14260 15534 14272
rect 15672 14260 15700 14288
rect 15528 14232 15700 14260
rect 15528 14220 15534 14232
rect 16206 14220 16212 14272
rect 16264 14260 16270 14272
rect 17788 14260 17816 14359
rect 16264 14232 17816 14260
rect 16264 14220 16270 14232
rect 1104 14170 18124 14192
rect 1104 14118 3737 14170
rect 3789 14118 3801 14170
rect 3853 14118 3865 14170
rect 3917 14118 3929 14170
rect 3981 14118 3993 14170
rect 4045 14118 7992 14170
rect 8044 14118 8056 14170
rect 8108 14118 8120 14170
rect 8172 14118 8184 14170
rect 8236 14118 8248 14170
rect 8300 14118 12247 14170
rect 12299 14118 12311 14170
rect 12363 14118 12375 14170
rect 12427 14118 12439 14170
rect 12491 14118 12503 14170
rect 12555 14118 16502 14170
rect 16554 14118 16566 14170
rect 16618 14118 16630 14170
rect 16682 14118 16694 14170
rect 16746 14118 16758 14170
rect 16810 14118 18124 14170
rect 1104 14096 18124 14118
rect 6365 14059 6423 14065
rect 6365 14025 6377 14059
rect 6411 14056 6423 14059
rect 6546 14056 6552 14068
rect 6411 14028 6552 14056
rect 6411 14025 6423 14028
rect 6365 14019 6423 14025
rect 6546 14016 6552 14028
rect 6604 14016 6610 14068
rect 7469 14059 7527 14065
rect 7469 14025 7481 14059
rect 7515 14056 7527 14059
rect 7650 14056 7656 14068
rect 7515 14028 7656 14056
rect 7515 14025 7527 14028
rect 7469 14019 7527 14025
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 7837 14059 7895 14065
rect 7837 14025 7849 14059
rect 7883 14056 7895 14059
rect 8386 14056 8392 14068
rect 7883 14028 8392 14056
rect 7883 14025 7895 14028
rect 7837 14019 7895 14025
rect 8386 14016 8392 14028
rect 8444 14016 8450 14068
rect 8496 14028 9076 14056
rect 2958 13948 2964 14000
rect 3016 13988 3022 14000
rect 4062 13988 4068 14000
rect 3016 13960 4068 13988
rect 3016 13948 3022 13960
rect 4062 13948 4068 13960
rect 4120 13988 4126 14000
rect 4341 13991 4399 13997
rect 4341 13988 4353 13991
rect 4120 13960 4353 13988
rect 4120 13948 4126 13960
rect 4341 13957 4353 13960
rect 4387 13957 4399 13991
rect 4341 13951 4399 13957
rect 4430 13948 4436 14000
rect 4488 13988 4494 14000
rect 6733 13991 6791 13997
rect 6733 13988 6745 13991
rect 4488 13960 6745 13988
rect 4488 13948 4494 13960
rect 6733 13957 6745 13960
rect 6779 13957 6791 13991
rect 7098 13988 7104 14000
rect 6733 13951 6791 13957
rect 6932 13960 7104 13988
rect 1946 13880 1952 13932
rect 2004 13880 2010 13932
rect 5166 13880 5172 13932
rect 5224 13920 5230 13932
rect 5261 13923 5319 13929
rect 5261 13920 5273 13923
rect 5224 13892 5273 13920
rect 5224 13880 5230 13892
rect 5261 13889 5273 13892
rect 5307 13889 5319 13923
rect 5261 13883 5319 13889
rect 6454 13880 6460 13932
rect 6512 13929 6518 13932
rect 6512 13923 6561 13929
rect 6512 13889 6515 13923
rect 6549 13889 6561 13923
rect 6512 13883 6561 13889
rect 6641 13923 6699 13929
rect 6641 13889 6653 13923
rect 6687 13889 6699 13923
rect 6641 13883 6699 13889
rect 6512 13880 6518 13883
rect 3329 13855 3387 13861
rect 3329 13821 3341 13855
rect 3375 13852 3387 13855
rect 3418 13852 3424 13864
rect 3375 13824 3424 13852
rect 3375 13821 3387 13824
rect 3329 13815 3387 13821
rect 3418 13812 3424 13824
rect 3476 13812 3482 13864
rect 5721 13855 5779 13861
rect 5721 13821 5733 13855
rect 5767 13852 5779 13855
rect 6656 13852 6684 13883
rect 6822 13880 6828 13932
rect 6880 13920 6886 13932
rect 6932 13929 6960 13960
rect 7098 13948 7104 13960
rect 7156 13988 7162 14000
rect 8496 13988 8524 14028
rect 7156 13960 8524 13988
rect 7156 13948 7162 13960
rect 8938 13948 8944 14000
rect 8996 13948 9002 14000
rect 6916 13923 6974 13929
rect 6916 13920 6928 13923
rect 6880 13892 6928 13920
rect 6880 13880 6886 13892
rect 6916 13889 6928 13892
rect 6962 13889 6974 13923
rect 6916 13883 6974 13889
rect 7009 13923 7067 13929
rect 7009 13889 7021 13923
rect 7055 13920 7067 13923
rect 7834 13920 7840 13932
rect 7055 13892 7840 13920
rect 7055 13889 7067 13892
rect 7009 13883 7067 13889
rect 7834 13880 7840 13892
rect 7892 13880 7898 13932
rect 7926 13880 7932 13932
rect 7984 13920 7990 13932
rect 9048 13920 9076 14028
rect 9306 14016 9312 14068
rect 9364 14016 9370 14068
rect 10042 14016 10048 14068
rect 10100 14016 10106 14068
rect 10134 14016 10140 14068
rect 10192 14016 10198 14068
rect 11146 14016 11152 14068
rect 11204 14056 11210 14068
rect 11609 14059 11667 14065
rect 11609 14056 11621 14059
rect 11204 14028 11621 14056
rect 11204 14016 11210 14028
rect 11609 14025 11621 14028
rect 11655 14025 11667 14059
rect 11609 14019 11667 14025
rect 11977 14059 12035 14065
rect 11977 14025 11989 14059
rect 12023 14056 12035 14059
rect 12618 14056 12624 14068
rect 12023 14028 12624 14056
rect 12023 14025 12035 14028
rect 11977 14019 12035 14025
rect 12618 14016 12624 14028
rect 12676 14016 12682 14068
rect 13538 14016 13544 14068
rect 13596 14056 13602 14068
rect 14737 14059 14795 14065
rect 14737 14056 14749 14059
rect 13596 14028 14749 14056
rect 13596 14016 13602 14028
rect 14737 14025 14749 14028
rect 14783 14025 14795 14059
rect 14737 14019 14795 14025
rect 15105 14059 15163 14065
rect 15105 14025 15117 14059
rect 15151 14056 15163 14059
rect 15933 14059 15991 14065
rect 15933 14056 15945 14059
rect 15151 14028 15945 14056
rect 15151 14025 15163 14028
rect 15105 14019 15163 14025
rect 15933 14025 15945 14028
rect 15979 14056 15991 14059
rect 16390 14056 16396 14068
rect 15979 14028 16396 14056
rect 15979 14025 15991 14028
rect 15933 14019 15991 14025
rect 16390 14016 16396 14028
rect 16448 14016 16454 14068
rect 16942 14016 16948 14068
rect 17000 14016 17006 14068
rect 12066 13948 12072 14000
rect 12124 13948 12130 14000
rect 12158 13948 12164 14000
rect 12216 13988 12222 14000
rect 12216 13960 14228 13988
rect 12216 13948 12222 13960
rect 9950 13920 9956 13932
rect 7984 13892 8892 13920
rect 9048 13892 9956 13920
rect 7984 13880 7990 13892
rect 8864 13861 8892 13892
rect 9950 13880 9956 13892
rect 10008 13880 10014 13932
rect 12618 13880 12624 13932
rect 12676 13880 12682 13932
rect 13188 13929 13216 13960
rect 13173 13923 13231 13929
rect 13173 13889 13185 13923
rect 13219 13889 13231 13923
rect 13173 13883 13231 13889
rect 13262 13880 13268 13932
rect 13320 13880 13326 13932
rect 13449 13923 13507 13929
rect 13449 13889 13461 13923
rect 13495 13920 13507 13923
rect 13906 13920 13912 13932
rect 13495 13892 13912 13920
rect 13495 13889 13507 13892
rect 13449 13883 13507 13889
rect 13906 13880 13912 13892
rect 13964 13880 13970 13932
rect 14200 13929 14228 13960
rect 15028 13960 15240 13988
rect 14185 13923 14243 13929
rect 14185 13889 14197 13923
rect 14231 13889 14243 13923
rect 14185 13883 14243 13889
rect 14274 13880 14280 13932
rect 14332 13880 14338 13932
rect 14458 13880 14464 13932
rect 14516 13880 14522 13932
rect 5767 13824 6684 13852
rect 8021 13855 8079 13861
rect 5767 13821 5779 13824
rect 5721 13815 5779 13821
rect 8021 13821 8033 13855
rect 8067 13821 8079 13855
rect 8021 13815 8079 13821
rect 8665 13855 8723 13861
rect 8665 13821 8677 13855
rect 8711 13821 8723 13855
rect 8665 13815 8723 13821
rect 8849 13855 8907 13861
rect 8849 13821 8861 13855
rect 8895 13852 8907 13855
rect 9858 13852 9864 13864
rect 8895 13824 9864 13852
rect 8895 13821 8907 13824
rect 8849 13815 8907 13821
rect 2958 13744 2964 13796
rect 3016 13784 3022 13796
rect 3016 13756 5672 13784
rect 3016 13744 3022 13756
rect 1670 13676 1676 13728
rect 1728 13716 1734 13728
rect 1765 13719 1823 13725
rect 1765 13716 1777 13719
rect 1728 13688 1777 13716
rect 1728 13676 1734 13688
rect 1765 13685 1777 13688
rect 1811 13685 1823 13719
rect 1765 13679 1823 13685
rect 2682 13676 2688 13728
rect 2740 13676 2746 13728
rect 5534 13676 5540 13728
rect 5592 13676 5598 13728
rect 5644 13716 5672 13756
rect 7650 13744 7656 13796
rect 7708 13784 7714 13796
rect 8036 13784 8064 13815
rect 7708 13756 8064 13784
rect 7708 13744 7714 13756
rect 8570 13744 8576 13796
rect 8628 13784 8634 13796
rect 8680 13784 8708 13815
rect 9858 13812 9864 13824
rect 9916 13812 9922 13864
rect 10321 13855 10379 13861
rect 10321 13821 10333 13855
rect 10367 13821 10379 13855
rect 10321 13815 10379 13821
rect 10336 13784 10364 13815
rect 10686 13812 10692 13864
rect 10744 13852 10750 13864
rect 11146 13852 11152 13864
rect 10744 13824 11152 13852
rect 10744 13812 10750 13824
rect 11146 13812 11152 13824
rect 11204 13852 11210 13864
rect 12161 13855 12219 13861
rect 12161 13852 12173 13855
rect 11204 13824 12173 13852
rect 11204 13812 11210 13824
rect 12161 13821 12173 13824
rect 12207 13821 12219 13855
rect 12161 13815 12219 13821
rect 13633 13787 13691 13793
rect 8628 13756 8708 13784
rect 8772 13756 13584 13784
rect 8628 13744 8634 13756
rect 8772 13716 8800 13756
rect 5644 13688 8800 13716
rect 9674 13676 9680 13728
rect 9732 13676 9738 13728
rect 12434 13676 12440 13728
rect 12492 13676 12498 13728
rect 13556 13716 13584 13756
rect 13633 13753 13645 13787
rect 13679 13784 13691 13787
rect 15028 13784 15056 13960
rect 15212 13920 15240 13960
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 16025 13991 16083 13997
rect 16025 13988 16037 13991
rect 15344 13960 16037 13988
rect 15344 13948 15350 13960
rect 16025 13957 16037 13960
rect 16071 13988 16083 13991
rect 16298 13988 16304 14000
rect 16071 13960 16304 13988
rect 16071 13957 16083 13960
rect 16025 13951 16083 13957
rect 16298 13948 16304 13960
rect 16356 13988 16362 14000
rect 16356 13960 17724 13988
rect 16356 13948 16362 13960
rect 17696 13929 17724 13960
rect 16761 13923 16819 13929
rect 15212 13892 15424 13920
rect 15194 13812 15200 13864
rect 15252 13812 15258 13864
rect 15289 13855 15347 13861
rect 15289 13821 15301 13855
rect 15335 13821 15347 13855
rect 15289 13815 15347 13821
rect 13679 13756 15056 13784
rect 13679 13753 13691 13756
rect 13633 13747 13691 13753
rect 15102 13744 15108 13796
rect 15160 13784 15166 13796
rect 15304 13784 15332 13815
rect 15160 13756 15332 13784
rect 15396 13784 15424 13892
rect 16761 13889 16773 13923
rect 16807 13889 16819 13923
rect 16761 13883 16819 13889
rect 17681 13923 17739 13929
rect 17681 13889 17693 13923
rect 17727 13889 17739 13923
rect 17681 13883 17739 13889
rect 15654 13812 15660 13864
rect 15712 13852 15718 13864
rect 16117 13855 16175 13861
rect 16117 13852 16129 13855
rect 15712 13824 16129 13852
rect 15712 13812 15718 13824
rect 16117 13821 16129 13824
rect 16163 13821 16175 13855
rect 16117 13815 16175 13821
rect 16776 13784 16804 13883
rect 15396 13756 16804 13784
rect 15160 13744 15166 13756
rect 14550 13716 14556 13728
rect 13556 13688 14556 13716
rect 14550 13676 14556 13688
rect 14608 13676 14614 13728
rect 14642 13676 14648 13728
rect 14700 13676 14706 13728
rect 15194 13676 15200 13728
rect 15252 13716 15258 13728
rect 15565 13719 15623 13725
rect 15565 13716 15577 13719
rect 15252 13688 15577 13716
rect 15252 13676 15258 13688
rect 15565 13685 15577 13688
rect 15611 13685 15623 13719
rect 15565 13679 15623 13685
rect 17126 13676 17132 13728
rect 17184 13676 17190 13728
rect 1104 13626 18124 13648
rect 1104 13574 3077 13626
rect 3129 13574 3141 13626
rect 3193 13574 3205 13626
rect 3257 13574 3269 13626
rect 3321 13574 3333 13626
rect 3385 13574 7332 13626
rect 7384 13574 7396 13626
rect 7448 13574 7460 13626
rect 7512 13574 7524 13626
rect 7576 13574 7588 13626
rect 7640 13574 11587 13626
rect 11639 13574 11651 13626
rect 11703 13574 11715 13626
rect 11767 13574 11779 13626
rect 11831 13574 11843 13626
rect 11895 13574 15842 13626
rect 15894 13574 15906 13626
rect 15958 13574 15970 13626
rect 16022 13574 16034 13626
rect 16086 13574 16098 13626
rect 16150 13574 18124 13626
rect 1104 13552 18124 13574
rect 3050 13472 3056 13524
rect 3108 13512 3114 13524
rect 10413 13515 10471 13521
rect 3108 13484 4384 13512
rect 3108 13472 3114 13484
rect 2777 13447 2835 13453
rect 2777 13413 2789 13447
rect 2823 13444 2835 13447
rect 2823 13416 3188 13444
rect 2823 13413 2835 13416
rect 2777 13407 2835 13413
rect 3050 13376 3056 13388
rect 2792 13348 3056 13376
rect 2792 13320 2820 13348
rect 3050 13336 3056 13348
rect 3108 13336 3114 13388
rect 3160 13385 3188 13416
rect 3145 13379 3203 13385
rect 3145 13345 3157 13379
rect 3191 13376 3203 13379
rect 3418 13376 3424 13388
rect 3191 13348 3424 13376
rect 3191 13345 3203 13348
rect 3145 13339 3203 13345
rect 3418 13336 3424 13348
rect 3476 13336 3482 13388
rect 4062 13336 4068 13388
rect 4120 13376 4126 13388
rect 4249 13379 4307 13385
rect 4249 13376 4261 13379
rect 4120 13348 4261 13376
rect 4120 13336 4126 13348
rect 4249 13345 4261 13348
rect 4295 13345 4307 13379
rect 4356 13376 4384 13484
rect 10413 13481 10425 13515
rect 10459 13512 10471 13515
rect 10502 13512 10508 13524
rect 10459 13484 10508 13512
rect 10459 13481 10471 13484
rect 10413 13475 10471 13481
rect 10502 13472 10508 13484
rect 10560 13472 10566 13524
rect 15562 13472 15568 13524
rect 15620 13512 15626 13524
rect 16025 13515 16083 13521
rect 16025 13512 16037 13515
rect 15620 13484 16037 13512
rect 15620 13472 15626 13484
rect 16025 13481 16037 13484
rect 16071 13512 16083 13515
rect 16206 13512 16212 13524
rect 16071 13484 16212 13512
rect 16071 13481 16083 13484
rect 16025 13475 16083 13481
rect 16206 13472 16212 13484
rect 16264 13472 16270 13524
rect 5718 13404 5724 13456
rect 5776 13444 5782 13456
rect 10134 13444 10140 13456
rect 5776 13416 10140 13444
rect 5776 13404 5782 13416
rect 10134 13404 10140 13416
rect 10192 13404 10198 13456
rect 10321 13447 10379 13453
rect 10321 13413 10333 13447
rect 10367 13413 10379 13447
rect 10321 13407 10379 13413
rect 12713 13447 12771 13453
rect 12713 13413 12725 13447
rect 12759 13413 12771 13447
rect 12713 13407 12771 13413
rect 9769 13379 9827 13385
rect 9769 13376 9781 13379
rect 4356 13348 9781 13376
rect 4249 13339 4307 13345
rect 9769 13345 9781 13348
rect 9815 13376 9827 13379
rect 10226 13376 10232 13388
rect 9815 13348 10232 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 10226 13336 10232 13348
rect 10284 13336 10290 13388
rect 10336 13376 10364 13407
rect 10336 13348 10824 13376
rect 1394 13268 1400 13320
rect 1452 13268 1458 13320
rect 1670 13317 1676 13320
rect 1664 13308 1676 13317
rect 1631 13280 1676 13308
rect 1664 13271 1676 13280
rect 1670 13268 1676 13271
rect 1728 13268 1734 13320
rect 2774 13268 2780 13320
rect 2832 13268 2838 13320
rect 3237 13311 3295 13317
rect 3237 13277 3249 13311
rect 3283 13308 3295 13311
rect 3510 13308 3516 13320
rect 3283 13280 3516 13308
rect 3283 13277 3295 13280
rect 3237 13271 3295 13277
rect 3510 13268 3516 13280
rect 3568 13268 3574 13320
rect 5994 13268 6000 13320
rect 6052 13268 6058 13320
rect 6546 13268 6552 13320
rect 6604 13268 6610 13320
rect 6730 13268 6736 13320
rect 6788 13308 6794 13320
rect 6825 13311 6883 13317
rect 6825 13308 6837 13311
rect 6788 13280 6837 13308
rect 6788 13268 6794 13280
rect 6825 13277 6837 13280
rect 6871 13277 6883 13311
rect 6825 13271 6883 13277
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13308 7067 13311
rect 7098 13308 7104 13320
rect 7055 13280 7104 13308
rect 7055 13277 7067 13280
rect 7009 13271 7067 13277
rect 7098 13268 7104 13280
rect 7156 13268 7162 13320
rect 9861 13311 9919 13317
rect 9861 13277 9873 13311
rect 9907 13308 9919 13311
rect 10318 13308 10324 13320
rect 9907 13280 10324 13308
rect 9907 13277 9919 13280
rect 9861 13271 9919 13277
rect 10318 13268 10324 13280
rect 10376 13268 10382 13320
rect 10594 13317 10600 13320
rect 10592 13308 10600 13317
rect 10555 13280 10600 13308
rect 10592 13271 10600 13280
rect 10594 13268 10600 13271
rect 10652 13268 10658 13320
rect 10686 13268 10692 13320
rect 10744 13268 10750 13320
rect 10796 13317 10824 13348
rect 10980 13348 11192 13376
rect 10980 13317 11008 13348
rect 10781 13311 10839 13317
rect 10781 13277 10793 13311
rect 10827 13277 10839 13311
rect 10964 13311 11022 13317
rect 10964 13308 10976 13311
rect 10781 13271 10839 13277
rect 10888 13280 10976 13308
rect 2590 13200 2596 13252
rect 2648 13240 2654 13252
rect 8570 13240 8576 13252
rect 2648 13212 8576 13240
rect 2648 13200 2654 13212
rect 8570 13200 8576 13212
rect 8628 13200 8634 13252
rect 9953 13243 10011 13249
rect 9953 13209 9965 13243
rect 9999 13240 10011 13243
rect 10042 13240 10048 13252
rect 9999 13212 10048 13240
rect 9999 13209 10011 13212
rect 9953 13203 10011 13209
rect 10042 13200 10048 13212
rect 10100 13200 10106 13252
rect 10134 13200 10140 13252
rect 10192 13240 10198 13252
rect 10888 13240 10916 13280
rect 10964 13277 10976 13280
rect 11010 13277 11022 13311
rect 10964 13271 11022 13277
rect 11057 13311 11115 13317
rect 11057 13277 11069 13311
rect 11103 13277 11115 13311
rect 11057 13271 11115 13277
rect 11072 13240 11100 13271
rect 10192 13212 10916 13240
rect 10980 13212 11100 13240
rect 11164 13240 11192 13348
rect 11330 13336 11336 13388
rect 11388 13336 11394 13388
rect 12728 13376 12756 13407
rect 14642 13404 14648 13456
rect 14700 13444 14706 13456
rect 17494 13444 17500 13456
rect 14700 13416 17500 13444
rect 14700 13404 14706 13416
rect 17494 13404 17500 13416
rect 17552 13404 17558 13456
rect 12986 13376 12992 13388
rect 12728 13348 12992 13376
rect 12986 13336 12992 13348
rect 13044 13376 13050 13388
rect 13357 13379 13415 13385
rect 13357 13376 13369 13379
rect 13044 13348 13369 13376
rect 13044 13336 13050 13348
rect 13357 13345 13369 13348
rect 13403 13345 13415 13379
rect 13357 13339 13415 13345
rect 16761 13379 16819 13385
rect 16761 13345 16773 13379
rect 16807 13376 16819 13379
rect 17218 13376 17224 13388
rect 16807 13348 17224 13376
rect 16807 13345 16819 13348
rect 16761 13339 16819 13345
rect 17218 13336 17224 13348
rect 17276 13336 17282 13388
rect 11600 13311 11658 13317
rect 11600 13277 11612 13311
rect 11646 13308 11658 13311
rect 12434 13308 12440 13320
rect 11646 13280 12440 13308
rect 11646 13277 11658 13280
rect 11600 13271 11658 13277
rect 12434 13268 12440 13280
rect 12492 13268 12498 13320
rect 12636 13280 13400 13308
rect 12636 13240 12664 13280
rect 13372 13252 13400 13280
rect 13814 13268 13820 13320
rect 13872 13308 13878 13320
rect 14737 13311 14795 13317
rect 14737 13308 14749 13311
rect 13872 13280 14749 13308
rect 13872 13268 13878 13280
rect 14737 13277 14749 13280
rect 14783 13277 14795 13311
rect 14737 13271 14795 13277
rect 15470 13268 15476 13320
rect 15528 13308 15534 13320
rect 16853 13311 16911 13317
rect 16853 13308 16865 13311
rect 15528 13280 16865 13308
rect 15528 13268 15534 13280
rect 16853 13277 16865 13280
rect 16899 13277 16911 13311
rect 16853 13271 16911 13277
rect 16945 13311 17003 13317
rect 16945 13277 16957 13311
rect 16991 13308 17003 13311
rect 17126 13308 17132 13320
rect 16991 13280 17132 13308
rect 16991 13277 17003 13280
rect 16945 13271 17003 13277
rect 13262 13240 13268 13252
rect 11164 13212 12664 13240
rect 12728 13212 13268 13240
rect 10192 13200 10198 13212
rect 3605 13175 3663 13181
rect 3605 13141 3617 13175
rect 3651 13172 3663 13175
rect 5810 13172 5816 13184
rect 3651 13144 5816 13172
rect 3651 13141 3663 13144
rect 3605 13135 3663 13141
rect 5810 13132 5816 13144
rect 5868 13132 5874 13184
rect 6362 13132 6368 13184
rect 6420 13132 6426 13184
rect 6638 13132 6644 13184
rect 6696 13172 6702 13184
rect 8938 13172 8944 13184
rect 6696 13144 8944 13172
rect 6696 13132 6702 13144
rect 8938 13132 8944 13144
rect 8996 13172 9002 13184
rect 10980 13172 11008 13212
rect 12728 13172 12756 13212
rect 13262 13200 13268 13212
rect 13320 13200 13326 13252
rect 13354 13200 13360 13252
rect 13412 13200 13418 13252
rect 14461 13243 14519 13249
rect 14461 13209 14473 13243
rect 14507 13240 14519 13243
rect 15562 13240 15568 13252
rect 14507 13212 15568 13240
rect 14507 13209 14519 13212
rect 14461 13203 14519 13209
rect 15562 13200 15568 13212
rect 15620 13200 15626 13252
rect 16868 13240 16896 13271
rect 17126 13268 17132 13280
rect 17184 13268 17190 13320
rect 17497 13311 17555 13317
rect 17497 13277 17509 13311
rect 17543 13277 17555 13311
rect 17497 13271 17555 13277
rect 17512 13240 17540 13271
rect 16868 13212 17540 13240
rect 17678 13200 17684 13252
rect 17736 13200 17742 13252
rect 8996 13144 12756 13172
rect 8996 13132 9002 13144
rect 12802 13132 12808 13184
rect 12860 13132 12866 13184
rect 14642 13132 14648 13184
rect 14700 13172 14706 13184
rect 15654 13172 15660 13184
rect 14700 13144 15660 13172
rect 14700 13132 14706 13144
rect 15654 13132 15660 13144
rect 15712 13132 15718 13184
rect 17313 13175 17371 13181
rect 17313 13141 17325 13175
rect 17359 13172 17371 13175
rect 17494 13172 17500 13184
rect 17359 13144 17500 13172
rect 17359 13141 17371 13144
rect 17313 13135 17371 13141
rect 17494 13132 17500 13144
rect 17552 13132 17558 13184
rect 1104 13082 18124 13104
rect 1104 13030 3737 13082
rect 3789 13030 3801 13082
rect 3853 13030 3865 13082
rect 3917 13030 3929 13082
rect 3981 13030 3993 13082
rect 4045 13030 7992 13082
rect 8044 13030 8056 13082
rect 8108 13030 8120 13082
rect 8172 13030 8184 13082
rect 8236 13030 8248 13082
rect 8300 13030 12247 13082
rect 12299 13030 12311 13082
rect 12363 13030 12375 13082
rect 12427 13030 12439 13082
rect 12491 13030 12503 13082
rect 12555 13030 16502 13082
rect 16554 13030 16566 13082
rect 16618 13030 16630 13082
rect 16682 13030 16694 13082
rect 16746 13030 16758 13082
rect 16810 13030 18124 13082
rect 1104 13008 18124 13030
rect 1946 12928 1952 12980
rect 2004 12968 2010 12980
rect 2133 12971 2191 12977
rect 2133 12968 2145 12971
rect 2004 12940 2145 12968
rect 2004 12928 2010 12940
rect 2133 12937 2145 12940
rect 2179 12937 2191 12971
rect 2133 12931 2191 12937
rect 2501 12971 2559 12977
rect 2501 12937 2513 12971
rect 2547 12968 2559 12971
rect 2682 12968 2688 12980
rect 2547 12940 2688 12968
rect 2547 12937 2559 12940
rect 2501 12931 2559 12937
rect 2682 12928 2688 12940
rect 2740 12928 2746 12980
rect 3237 12971 3295 12977
rect 3237 12937 3249 12971
rect 3283 12968 3295 12971
rect 3418 12968 3424 12980
rect 3283 12940 3424 12968
rect 3283 12937 3295 12940
rect 3237 12931 3295 12937
rect 3418 12928 3424 12940
rect 3476 12928 3482 12980
rect 5169 12971 5227 12977
rect 3620 12940 5120 12968
rect 1026 12860 1032 12912
rect 1084 12900 1090 12912
rect 1489 12903 1547 12909
rect 1489 12900 1501 12903
rect 1084 12872 1501 12900
rect 1084 12860 1090 12872
rect 1489 12869 1501 12872
rect 1535 12869 1547 12903
rect 1489 12863 1547 12869
rect 3329 12903 3387 12909
rect 3329 12869 3341 12903
rect 3375 12900 3387 12903
rect 3510 12900 3516 12912
rect 3375 12872 3516 12900
rect 3375 12869 3387 12872
rect 3329 12863 3387 12869
rect 3510 12860 3516 12872
rect 3568 12860 3574 12912
rect 2498 12724 2504 12776
rect 2556 12764 2562 12776
rect 2593 12767 2651 12773
rect 2593 12764 2605 12767
rect 2556 12736 2605 12764
rect 2556 12724 2562 12736
rect 2593 12733 2605 12736
rect 2639 12733 2651 12767
rect 2593 12727 2651 12733
rect 2682 12724 2688 12776
rect 2740 12724 2746 12776
rect 2958 12724 2964 12776
rect 3016 12764 3022 12776
rect 3053 12767 3111 12773
rect 3053 12764 3065 12767
rect 3016 12736 3065 12764
rect 3016 12724 3022 12736
rect 3053 12733 3065 12736
rect 3099 12733 3111 12767
rect 3053 12727 3111 12733
rect 1394 12656 1400 12708
rect 1452 12696 1458 12708
rect 2866 12696 2872 12708
rect 1452 12668 2872 12696
rect 1452 12656 1458 12668
rect 2866 12656 2872 12668
rect 2924 12656 2930 12708
rect 1765 12631 1823 12637
rect 1765 12597 1777 12631
rect 1811 12628 1823 12631
rect 3620 12628 3648 12940
rect 3694 12792 3700 12844
rect 3752 12832 3758 12844
rect 3789 12835 3847 12841
rect 3789 12832 3801 12835
rect 3752 12804 3801 12832
rect 3752 12792 3758 12804
rect 3789 12801 3801 12804
rect 3835 12832 3847 12835
rect 3878 12832 3884 12844
rect 3835 12804 3884 12832
rect 3835 12801 3847 12804
rect 3789 12795 3847 12801
rect 3878 12792 3884 12804
rect 3936 12792 3942 12844
rect 4062 12841 4068 12844
rect 4056 12795 4068 12841
rect 4062 12792 4068 12795
rect 4120 12792 4126 12844
rect 5092 12832 5120 12940
rect 5169 12937 5181 12971
rect 5215 12968 5227 12971
rect 5534 12968 5540 12980
rect 5215 12940 5540 12968
rect 5215 12937 5227 12940
rect 5169 12931 5227 12937
rect 5534 12928 5540 12940
rect 5592 12928 5598 12980
rect 6181 12971 6239 12977
rect 6181 12937 6193 12971
rect 6227 12968 6239 12971
rect 6270 12968 6276 12980
rect 6227 12940 6276 12968
rect 6227 12937 6239 12940
rect 6181 12931 6239 12937
rect 6270 12928 6276 12940
rect 6328 12928 6334 12980
rect 6825 12971 6883 12977
rect 6825 12937 6837 12971
rect 6871 12937 6883 12971
rect 6825 12931 6883 12937
rect 9232 12940 10180 12968
rect 5810 12860 5816 12912
rect 5868 12860 5874 12912
rect 6840 12900 6868 12931
rect 7162 12903 7220 12909
rect 7162 12900 7174 12903
rect 6840 12872 7174 12900
rect 7162 12869 7174 12872
rect 7208 12869 7220 12903
rect 7162 12863 7220 12869
rect 9232 12844 9260 12940
rect 9674 12860 9680 12912
rect 9732 12900 9738 12912
rect 10045 12903 10103 12909
rect 10045 12900 10057 12903
rect 9732 12872 10057 12900
rect 9732 12860 9738 12872
rect 10045 12869 10057 12872
rect 10091 12869 10103 12903
rect 10152 12900 10180 12940
rect 10410 12928 10416 12980
rect 10468 12928 10474 12980
rect 12066 12928 12072 12980
rect 12124 12968 12130 12980
rect 12161 12971 12219 12977
rect 12161 12968 12173 12971
rect 12124 12940 12173 12968
rect 12124 12928 12130 12940
rect 12161 12937 12173 12940
rect 12207 12937 12219 12971
rect 12161 12931 12219 12937
rect 12618 12928 12624 12980
rect 12676 12928 12682 12980
rect 13909 12971 13967 12977
rect 13909 12937 13921 12971
rect 13955 12968 13967 12971
rect 14366 12968 14372 12980
rect 13955 12940 14372 12968
rect 13955 12937 13967 12940
rect 13909 12931 13967 12937
rect 14366 12928 14372 12940
rect 14424 12928 14430 12980
rect 14458 12928 14464 12980
rect 14516 12968 14522 12980
rect 14645 12971 14703 12977
rect 14645 12968 14657 12971
rect 14516 12940 14657 12968
rect 14516 12928 14522 12940
rect 14645 12937 14657 12940
rect 14691 12937 14703 12971
rect 14645 12931 14703 12937
rect 17405 12971 17463 12977
rect 17405 12937 17417 12971
rect 17451 12937 17463 12971
rect 17405 12931 17463 12937
rect 12253 12903 12311 12909
rect 10152 12872 11376 12900
rect 10045 12863 10103 12869
rect 5718 12841 5724 12844
rect 5537 12835 5595 12841
rect 5537 12832 5549 12835
rect 5092 12804 5549 12832
rect 5537 12801 5549 12804
rect 5583 12801 5595 12835
rect 5537 12795 5595 12801
rect 5685 12835 5724 12841
rect 5685 12801 5697 12835
rect 5685 12795 5724 12801
rect 5552 12696 5580 12795
rect 5718 12792 5724 12795
rect 5776 12792 5782 12844
rect 5902 12792 5908 12844
rect 5960 12792 5966 12844
rect 6043 12835 6101 12841
rect 6043 12801 6055 12835
rect 6089 12832 6101 12835
rect 6362 12832 6368 12844
rect 6089 12804 6368 12832
rect 6089 12801 6101 12804
rect 6043 12795 6101 12801
rect 6362 12792 6368 12804
rect 6420 12792 6426 12844
rect 6641 12835 6699 12841
rect 6641 12801 6653 12835
rect 6687 12832 6699 12835
rect 7006 12832 7012 12844
rect 6687 12804 7012 12832
rect 6687 12801 6699 12804
rect 6641 12795 6699 12801
rect 7006 12792 7012 12804
rect 7064 12792 7070 12844
rect 9214 12792 9220 12844
rect 9272 12792 9278 12844
rect 9950 12841 9956 12844
rect 9769 12835 9827 12841
rect 9769 12832 9781 12835
rect 9600 12804 9781 12832
rect 6914 12724 6920 12776
rect 6972 12724 6978 12776
rect 8941 12767 8999 12773
rect 8941 12764 8953 12767
rect 8312 12736 8953 12764
rect 5626 12696 5632 12708
rect 5552 12668 5632 12696
rect 5626 12656 5632 12668
rect 5684 12696 5690 12708
rect 6638 12696 6644 12708
rect 5684 12668 6644 12696
rect 5684 12656 5690 12668
rect 6638 12656 6644 12668
rect 6696 12656 6702 12708
rect 1811 12600 3648 12628
rect 3697 12631 3755 12637
rect 1811 12597 1823 12600
rect 1765 12591 1823 12597
rect 3697 12597 3709 12631
rect 3743 12628 3755 12631
rect 4430 12628 4436 12640
rect 3743 12600 4436 12628
rect 3743 12597 3755 12600
rect 3697 12591 3755 12597
rect 4430 12588 4436 12600
rect 4488 12588 4494 12640
rect 7098 12588 7104 12640
rect 7156 12628 7162 12640
rect 8312 12637 8340 12736
rect 8941 12733 8953 12736
rect 8987 12733 8999 12767
rect 8941 12727 8999 12733
rect 9600 12696 9628 12804
rect 9769 12801 9781 12804
rect 9815 12801 9827 12835
rect 9769 12795 9827 12801
rect 9917 12835 9956 12841
rect 9917 12801 9929 12835
rect 9917 12795 9956 12801
rect 9950 12792 9956 12795
rect 10008 12792 10014 12844
rect 10137 12835 10195 12841
rect 10137 12801 10149 12835
rect 10183 12801 10195 12835
rect 10137 12795 10195 12801
rect 10275 12835 10333 12841
rect 10275 12801 10287 12835
rect 10321 12832 10333 12835
rect 10689 12835 10747 12841
rect 10689 12832 10701 12835
rect 10321 12804 10701 12832
rect 10321 12801 10333 12804
rect 10275 12795 10333 12801
rect 10689 12801 10701 12804
rect 10735 12801 10747 12835
rect 10689 12795 10747 12801
rect 9677 12767 9735 12773
rect 9677 12733 9689 12767
rect 9723 12764 9735 12767
rect 10152 12764 10180 12795
rect 10870 12792 10876 12844
rect 10928 12792 10934 12844
rect 11149 12835 11207 12841
rect 11149 12801 11161 12835
rect 11195 12832 11207 12835
rect 11238 12832 11244 12844
rect 11195 12804 11244 12832
rect 11195 12801 11207 12804
rect 11149 12795 11207 12801
rect 11238 12792 11244 12804
rect 11296 12792 11302 12844
rect 11348 12841 11376 12872
rect 12253 12869 12265 12903
rect 12299 12900 12311 12903
rect 12802 12900 12808 12912
rect 12299 12872 12808 12900
rect 12299 12869 12311 12872
rect 12253 12863 12311 12869
rect 12802 12860 12808 12872
rect 12860 12860 12866 12912
rect 13538 12860 13544 12912
rect 13596 12860 13602 12912
rect 14277 12903 14335 12909
rect 14277 12869 14289 12903
rect 14323 12900 14335 12903
rect 15194 12900 15200 12912
rect 14323 12872 15200 12900
rect 14323 12869 14335 12872
rect 14277 12863 14335 12869
rect 15194 12860 15200 12872
rect 15252 12860 15258 12912
rect 16240 12903 16298 12909
rect 16240 12869 16252 12903
rect 16286 12900 16298 12903
rect 17420 12900 17448 12931
rect 16286 12872 17448 12900
rect 16286 12869 16298 12872
rect 16240 12863 16298 12869
rect 11333 12835 11391 12841
rect 11333 12801 11345 12835
rect 11379 12832 11391 12835
rect 12434 12832 12440 12844
rect 11379 12804 12440 12832
rect 11379 12801 11391 12804
rect 11333 12795 11391 12801
rect 12434 12792 12440 12804
rect 12492 12792 12498 12844
rect 12710 12792 12716 12844
rect 12768 12792 12774 12844
rect 13262 12792 13268 12844
rect 13320 12792 13326 12844
rect 13354 12792 13360 12844
rect 13412 12832 13418 12844
rect 13633 12835 13691 12841
rect 13412 12804 13457 12832
rect 13412 12792 13418 12804
rect 13633 12801 13645 12835
rect 13679 12801 13691 12835
rect 13633 12795 13691 12801
rect 9723 12736 10180 12764
rect 9723 12733 9735 12736
rect 9677 12727 9735 12733
rect 12066 12724 12072 12776
rect 12124 12724 12130 12776
rect 13173 12767 13231 12773
rect 13173 12733 13185 12767
rect 13219 12764 13231 12767
rect 13648 12764 13676 12795
rect 13722 12792 13728 12844
rect 13780 12841 13786 12844
rect 14182 12841 14188 12844
rect 13780 12832 13788 12841
rect 14001 12835 14059 12841
rect 13780 12804 13825 12832
rect 13780 12795 13788 12804
rect 14001 12801 14013 12835
rect 14047 12801 14059 12835
rect 14001 12795 14059 12801
rect 14149 12835 14188 12841
rect 14149 12801 14161 12835
rect 14149 12795 14188 12801
rect 13780 12792 13786 12795
rect 13219 12736 13676 12764
rect 14016 12764 14044 12795
rect 14182 12792 14188 12795
rect 14240 12792 14246 12844
rect 14366 12792 14372 12844
rect 14424 12792 14430 12844
rect 14458 12792 14464 12844
rect 14516 12841 14522 12844
rect 14516 12832 14524 12841
rect 14516 12804 14561 12832
rect 14516 12795 14524 12804
rect 14516 12792 14522 12795
rect 16574 12792 16580 12844
rect 16632 12832 16638 12844
rect 17589 12835 17647 12841
rect 17589 12832 17601 12835
rect 16632 12804 17601 12832
rect 16632 12792 16638 12804
rect 17589 12801 17601 12804
rect 17635 12801 17647 12835
rect 17589 12795 17647 12801
rect 14550 12764 14556 12776
rect 14016 12736 14556 12764
rect 13219 12733 13231 12736
rect 13173 12727 13231 12733
rect 14016 12696 14044 12736
rect 14550 12724 14556 12736
rect 14608 12724 14614 12776
rect 16482 12724 16488 12776
rect 16540 12724 16546 12776
rect 17221 12767 17279 12773
rect 17221 12733 17233 12767
rect 17267 12733 17279 12767
rect 17221 12727 17279 12733
rect 17236 12696 17264 12727
rect 9600 12668 14044 12696
rect 16500 12668 17264 12696
rect 9692 12640 9720 12668
rect 8297 12631 8355 12637
rect 8297 12628 8309 12631
rect 7156 12600 8309 12628
rect 7156 12588 7162 12600
rect 8297 12597 8309 12600
rect 8343 12597 8355 12631
rect 8297 12591 8355 12597
rect 8386 12588 8392 12640
rect 8444 12588 8450 12640
rect 9398 12588 9404 12640
rect 9456 12588 9462 12640
rect 9674 12588 9680 12640
rect 9732 12588 9738 12640
rect 10226 12588 10232 12640
rect 10284 12628 10290 12640
rect 12618 12628 12624 12640
rect 10284 12600 12624 12628
rect 10284 12588 10290 12600
rect 12618 12588 12624 12600
rect 12676 12588 12682 12640
rect 12986 12588 12992 12640
rect 13044 12588 13050 12640
rect 14918 12588 14924 12640
rect 14976 12628 14982 12640
rect 15105 12631 15163 12637
rect 15105 12628 15117 12631
rect 14976 12600 15117 12628
rect 14976 12588 14982 12600
rect 15105 12597 15117 12600
rect 15151 12628 15163 12631
rect 16500 12628 16528 12668
rect 15151 12600 16528 12628
rect 15151 12597 15163 12600
rect 15105 12591 15163 12597
rect 16666 12588 16672 12640
rect 16724 12588 16730 12640
rect 1104 12538 18124 12560
rect 1104 12486 3077 12538
rect 3129 12486 3141 12538
rect 3193 12486 3205 12538
rect 3257 12486 3269 12538
rect 3321 12486 3333 12538
rect 3385 12486 7332 12538
rect 7384 12486 7396 12538
rect 7448 12486 7460 12538
rect 7512 12486 7524 12538
rect 7576 12486 7588 12538
rect 7640 12486 11587 12538
rect 11639 12486 11651 12538
rect 11703 12486 11715 12538
rect 11767 12486 11779 12538
rect 11831 12486 11843 12538
rect 11895 12486 15842 12538
rect 15894 12486 15906 12538
rect 15958 12486 15970 12538
rect 16022 12486 16034 12538
rect 16086 12486 16098 12538
rect 16150 12486 18124 12538
rect 1104 12464 18124 12486
rect 3973 12427 4031 12433
rect 3973 12393 3985 12427
rect 4019 12424 4031 12427
rect 4062 12424 4068 12436
rect 4019 12396 4068 12424
rect 4019 12393 4031 12396
rect 3973 12387 4031 12393
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 5813 12427 5871 12433
rect 5813 12393 5825 12427
rect 5859 12424 5871 12427
rect 5902 12424 5908 12436
rect 5859 12396 5908 12424
rect 5859 12393 5871 12396
rect 5813 12387 5871 12393
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 5997 12427 6055 12433
rect 5997 12393 6009 12427
rect 6043 12393 6055 12427
rect 5997 12387 6055 12393
rect 6365 12427 6423 12433
rect 6365 12393 6377 12427
rect 6411 12424 6423 12427
rect 6454 12424 6460 12436
rect 6411 12396 6460 12424
rect 6411 12393 6423 12396
rect 6365 12387 6423 12393
rect 2498 12248 2504 12300
rect 2556 12288 2562 12300
rect 2556 12260 4568 12288
rect 2556 12248 2562 12260
rect 1302 12180 1308 12232
rect 1360 12220 1366 12232
rect 1489 12223 1547 12229
rect 1489 12220 1501 12223
rect 1360 12192 1501 12220
rect 1360 12180 1366 12192
rect 1489 12189 1501 12192
rect 1535 12189 1547 12223
rect 1489 12183 1547 12189
rect 2038 12180 2044 12232
rect 2096 12220 2102 12232
rect 2133 12223 2191 12229
rect 2133 12220 2145 12223
rect 2096 12192 2145 12220
rect 2096 12180 2102 12192
rect 2133 12189 2145 12192
rect 2179 12189 2191 12223
rect 2133 12183 2191 12189
rect 2866 12180 2872 12232
rect 2924 12220 2930 12232
rect 3329 12223 3387 12229
rect 3329 12220 3341 12223
rect 2924 12192 3341 12220
rect 2924 12180 2930 12192
rect 3329 12189 3341 12192
rect 3375 12189 3387 12223
rect 3329 12183 3387 12189
rect 4157 12223 4215 12229
rect 4157 12189 4169 12223
rect 4203 12220 4215 12223
rect 4203 12192 4292 12220
rect 4203 12189 4215 12192
rect 4157 12183 4215 12189
rect 1762 12044 1768 12096
rect 1820 12044 1826 12096
rect 1854 12044 1860 12096
rect 1912 12084 1918 12096
rect 1949 12087 2007 12093
rect 1949 12084 1961 12087
rect 1912 12056 1961 12084
rect 1912 12044 1918 12056
rect 1949 12053 1961 12056
rect 1995 12053 2007 12087
rect 1949 12047 2007 12053
rect 2406 12044 2412 12096
rect 2464 12084 2470 12096
rect 4264 12093 4292 12192
rect 2777 12087 2835 12093
rect 2777 12084 2789 12087
rect 2464 12056 2789 12084
rect 2464 12044 2470 12056
rect 2777 12053 2789 12056
rect 2823 12053 2835 12087
rect 2777 12047 2835 12053
rect 4249 12087 4307 12093
rect 4249 12053 4261 12087
rect 4295 12053 4307 12087
rect 4540 12084 4568 12260
rect 4798 12248 4804 12300
rect 4856 12248 4862 12300
rect 5534 12248 5540 12300
rect 5592 12288 5598 12300
rect 5721 12291 5779 12297
rect 5721 12288 5733 12291
rect 5592 12260 5733 12288
rect 5592 12248 5598 12260
rect 5721 12257 5733 12260
rect 5767 12288 5779 12291
rect 6012 12288 6040 12387
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7101 12427 7159 12433
rect 7101 12424 7113 12427
rect 7064 12396 7113 12424
rect 7064 12384 7070 12396
rect 7101 12393 7113 12396
rect 7147 12393 7159 12427
rect 7834 12424 7840 12436
rect 7101 12387 7159 12393
rect 7484 12396 7840 12424
rect 6086 12316 6092 12368
rect 6144 12356 6150 12368
rect 7484 12356 7512 12396
rect 7834 12384 7840 12396
rect 7892 12424 7898 12436
rect 8202 12424 8208 12436
rect 7892 12396 8208 12424
rect 7892 12384 7898 12396
rect 8202 12384 8208 12396
rect 8260 12424 8266 12436
rect 8260 12396 9343 12424
rect 8260 12384 8266 12396
rect 8386 12356 8392 12368
rect 6144 12328 7512 12356
rect 7576 12328 8392 12356
rect 6144 12316 6150 12328
rect 5767 12260 6040 12288
rect 5767 12257 5779 12260
rect 5721 12251 5779 12257
rect 6730 12248 6736 12300
rect 6788 12288 6794 12300
rect 7576 12297 7604 12328
rect 8386 12316 8392 12328
rect 8444 12316 8450 12368
rect 9315 12356 9343 12396
rect 9398 12384 9404 12436
rect 9456 12424 9462 12436
rect 9493 12427 9551 12433
rect 9493 12424 9505 12427
rect 9456 12396 9505 12424
rect 9456 12384 9462 12396
rect 9493 12393 9505 12396
rect 9539 12393 9551 12427
rect 9493 12387 9551 12393
rect 10594 12384 10600 12436
rect 10652 12424 10658 12436
rect 10689 12427 10747 12433
rect 10689 12424 10701 12427
rect 10652 12396 10701 12424
rect 10652 12384 10658 12396
rect 10689 12393 10701 12396
rect 10735 12393 10747 12427
rect 10689 12387 10747 12393
rect 12986 12384 12992 12436
rect 13044 12384 13050 12436
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 14277 12427 14335 12433
rect 14277 12424 14289 12427
rect 13780 12396 14289 12424
rect 13780 12384 13786 12396
rect 14277 12393 14289 12396
rect 14323 12393 14335 12427
rect 14277 12387 14335 12393
rect 16298 12384 16304 12436
rect 16356 12384 16362 12436
rect 16390 12384 16396 12436
rect 16448 12384 16454 12436
rect 9674 12356 9680 12368
rect 9315 12328 9680 12356
rect 9674 12316 9680 12328
rect 9732 12316 9738 12368
rect 13265 12359 13323 12365
rect 13265 12325 13277 12359
rect 13311 12356 13323 12359
rect 14366 12356 14372 12368
rect 13311 12328 14372 12356
rect 13311 12325 13323 12328
rect 13265 12319 13323 12325
rect 14366 12316 14372 12328
rect 14424 12316 14430 12368
rect 7561 12291 7619 12297
rect 6788 12260 7512 12288
rect 6788 12248 6794 12260
rect 5166 12180 5172 12232
rect 5224 12220 5230 12232
rect 5442 12220 5448 12232
rect 5224 12192 5448 12220
rect 5224 12180 5230 12192
rect 5442 12180 5448 12192
rect 5500 12220 5506 12232
rect 6273 12223 6331 12229
rect 6273 12220 6285 12223
rect 5500 12192 6285 12220
rect 5500 12180 5506 12192
rect 6273 12189 6285 12192
rect 6319 12189 6331 12223
rect 6273 12183 6331 12189
rect 6546 12180 6552 12232
rect 6604 12180 6610 12232
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12189 6883 12223
rect 6825 12183 6883 12189
rect 7009 12223 7067 12229
rect 7009 12189 7021 12223
rect 7055 12220 7067 12223
rect 7098 12220 7104 12232
rect 7055 12192 7104 12220
rect 7055 12189 7067 12192
rect 7009 12183 7067 12189
rect 4617 12155 4675 12161
rect 4617 12121 4629 12155
rect 4663 12152 4675 12155
rect 5077 12155 5135 12161
rect 5077 12152 5089 12155
rect 4663 12124 5089 12152
rect 4663 12121 4675 12124
rect 4617 12115 4675 12121
rect 5077 12121 5089 12124
rect 5123 12121 5135 12155
rect 6840 12152 6868 12183
rect 7098 12180 7104 12192
rect 7156 12180 7162 12232
rect 7484 12220 7512 12260
rect 7561 12257 7573 12291
rect 7607 12257 7619 12291
rect 7561 12251 7619 12257
rect 7745 12291 7803 12297
rect 7745 12257 7757 12291
rect 7791 12288 7803 12291
rect 7834 12288 7840 12300
rect 7791 12260 7840 12288
rect 7791 12257 7803 12260
rect 7745 12251 7803 12257
rect 7834 12248 7840 12260
rect 7892 12248 7898 12300
rect 9861 12291 9919 12297
rect 8312 12260 9444 12288
rect 8312 12220 8340 12260
rect 7484 12192 8340 12220
rect 8386 12180 8392 12232
rect 8444 12180 8450 12232
rect 8938 12180 8944 12232
rect 8996 12180 9002 12232
rect 9416 12229 9444 12260
rect 9861 12257 9873 12291
rect 9907 12288 9919 12291
rect 10686 12288 10692 12300
rect 9907 12260 10692 12288
rect 9907 12257 9919 12260
rect 9861 12251 9919 12257
rect 10686 12248 10692 12260
rect 10744 12248 10750 12300
rect 15102 12288 15108 12300
rect 10888 12260 13860 12288
rect 10888 12229 10916 12260
rect 13832 12232 13860 12260
rect 14844 12260 15108 12288
rect 14844 12232 14872 12260
rect 15102 12248 15108 12260
rect 15160 12248 15166 12300
rect 15194 12248 15200 12300
rect 15252 12288 15258 12300
rect 15657 12291 15715 12297
rect 15657 12288 15669 12291
rect 15252 12260 15669 12288
rect 15252 12248 15258 12260
rect 15657 12257 15669 12260
rect 15703 12257 15715 12291
rect 15657 12251 15715 12257
rect 15841 12291 15899 12297
rect 15841 12257 15853 12291
rect 15887 12288 15899 12291
rect 16666 12288 16672 12300
rect 15887 12260 16672 12288
rect 15887 12257 15899 12260
rect 15841 12251 15899 12257
rect 16666 12248 16672 12260
rect 16724 12248 16730 12300
rect 9401 12223 9459 12229
rect 9401 12189 9413 12223
rect 9447 12189 9459 12223
rect 9401 12183 9459 12189
rect 10873 12223 10931 12229
rect 10873 12189 10885 12223
rect 10919 12189 10931 12223
rect 10873 12183 10931 12189
rect 11149 12223 11207 12229
rect 11149 12189 11161 12223
rect 11195 12189 11207 12223
rect 11149 12183 11207 12189
rect 7190 12152 7196 12164
rect 6840 12124 7196 12152
rect 5077 12115 5135 12121
rect 7190 12112 7196 12124
rect 7248 12152 7254 12164
rect 9214 12152 9220 12164
rect 7248 12124 9220 12152
rect 7248 12112 7254 12124
rect 9214 12112 9220 12124
rect 9272 12112 9278 12164
rect 9416 12152 9444 12183
rect 11164 12152 11192 12183
rect 11238 12180 11244 12232
rect 11296 12220 11302 12232
rect 11333 12223 11391 12229
rect 11333 12220 11345 12223
rect 11296 12192 11345 12220
rect 11296 12180 11302 12192
rect 11333 12189 11345 12192
rect 11379 12189 11391 12223
rect 11333 12183 11391 12189
rect 12434 12180 12440 12232
rect 12492 12220 12498 12232
rect 12802 12220 12808 12232
rect 12492 12192 12808 12220
rect 12492 12180 12498 12192
rect 12802 12180 12808 12192
rect 12860 12180 12866 12232
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 14461 12223 14519 12229
rect 14461 12220 14473 12223
rect 13872 12192 14473 12220
rect 13872 12180 13878 12192
rect 14461 12189 14473 12192
rect 14507 12189 14519 12223
rect 14461 12183 14519 12189
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 14826 12220 14832 12232
rect 14783 12192 14832 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 12710 12152 12716 12164
rect 9416 12124 12716 12152
rect 12710 12112 12716 12124
rect 12768 12112 12774 12164
rect 4709 12087 4767 12093
rect 4709 12084 4721 12087
rect 4540 12056 4721 12084
rect 4249 12047 4307 12053
rect 4709 12053 4721 12056
rect 4755 12084 4767 12087
rect 7469 12087 7527 12093
rect 7469 12084 7481 12087
rect 4755 12056 7481 12084
rect 4755 12053 4767 12056
rect 4709 12047 4767 12053
rect 7469 12053 7481 12056
rect 7515 12053 7527 12087
rect 7469 12047 7527 12053
rect 8481 12087 8539 12093
rect 8481 12053 8493 12087
rect 8527 12084 8539 12087
rect 8570 12084 8576 12096
rect 8527 12056 8576 12084
rect 8527 12053 8539 12056
rect 8481 12047 8539 12053
rect 8570 12044 8576 12056
rect 8628 12044 8634 12096
rect 9030 12044 9036 12096
rect 9088 12044 9094 12096
rect 12618 12044 12624 12096
rect 12676 12084 12682 12096
rect 13998 12084 14004 12096
rect 12676 12056 14004 12084
rect 12676 12044 12682 12056
rect 13998 12044 14004 12056
rect 14056 12084 14062 12096
rect 14752 12084 14780 12183
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 14918 12180 14924 12232
rect 14976 12180 14982 12232
rect 16390 12180 16396 12232
rect 16448 12220 16454 12232
rect 17773 12223 17831 12229
rect 17773 12220 17785 12223
rect 16448 12192 17785 12220
rect 16448 12180 16454 12192
rect 17773 12189 17785 12192
rect 17819 12189 17831 12223
rect 17773 12183 17831 12189
rect 15654 12112 15660 12164
rect 15712 12152 15718 12164
rect 15933 12155 15991 12161
rect 15933 12152 15945 12155
rect 15712 12124 15945 12152
rect 15712 12112 15718 12124
rect 15933 12121 15945 12124
rect 15979 12121 15991 12155
rect 15933 12115 15991 12121
rect 17528 12155 17586 12161
rect 17528 12121 17540 12155
rect 17574 12152 17586 12155
rect 17678 12152 17684 12164
rect 17574 12124 17684 12152
rect 17574 12121 17586 12124
rect 17528 12115 17586 12121
rect 17678 12112 17684 12124
rect 17736 12112 17742 12164
rect 14056 12056 14780 12084
rect 14056 12044 14062 12056
rect 1104 11994 18124 12016
rect 1104 11942 3737 11994
rect 3789 11942 3801 11994
rect 3853 11942 3865 11994
rect 3917 11942 3929 11994
rect 3981 11942 3993 11994
rect 4045 11942 7992 11994
rect 8044 11942 8056 11994
rect 8108 11942 8120 11994
rect 8172 11942 8184 11994
rect 8236 11942 8248 11994
rect 8300 11942 12247 11994
rect 12299 11942 12311 11994
rect 12363 11942 12375 11994
rect 12427 11942 12439 11994
rect 12491 11942 12503 11994
rect 12555 11942 16502 11994
rect 16554 11942 16566 11994
rect 16618 11942 16630 11994
rect 16682 11942 16694 11994
rect 16746 11942 16758 11994
rect 16810 11942 18124 11994
rect 1104 11920 18124 11942
rect 4798 11840 4804 11892
rect 4856 11880 4862 11892
rect 8662 11880 8668 11892
rect 4856 11852 8668 11880
rect 4856 11840 4862 11852
rect 8662 11840 8668 11852
rect 8720 11840 8726 11892
rect 8757 11883 8815 11889
rect 8757 11849 8769 11883
rect 8803 11849 8815 11883
rect 13998 11880 14004 11892
rect 8757 11843 8815 11849
rect 13832 11852 14004 11880
rect 1762 11772 1768 11824
rect 1820 11812 1826 11824
rect 5534 11812 5540 11824
rect 1820 11784 5540 11812
rect 1820 11772 1826 11784
rect 5534 11772 5540 11784
rect 5592 11772 5598 11824
rect 1854 11753 1860 11756
rect 1848 11744 1860 11753
rect 1815 11716 1860 11744
rect 1848 11707 1860 11716
rect 1854 11704 1860 11707
rect 1912 11704 1918 11756
rect 3602 11704 3608 11756
rect 3660 11704 3666 11756
rect 3878 11753 3884 11756
rect 3872 11707 3884 11753
rect 3878 11704 3884 11707
rect 3936 11704 3942 11756
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11744 6607 11747
rect 6638 11744 6644 11756
rect 6595 11716 6644 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 6638 11704 6644 11716
rect 6696 11704 6702 11756
rect 6730 11704 6736 11756
rect 6788 11744 6794 11756
rect 6825 11747 6883 11753
rect 6825 11744 6837 11747
rect 6788 11716 6837 11744
rect 6788 11704 6794 11716
rect 6825 11713 6837 11716
rect 6871 11713 6883 11747
rect 6825 11707 6883 11713
rect 7006 11704 7012 11756
rect 7064 11704 7070 11756
rect 8665 11747 8723 11753
rect 8665 11713 8677 11747
rect 8711 11744 8723 11747
rect 8772 11744 8800 11843
rect 9217 11815 9275 11821
rect 9217 11781 9229 11815
rect 9263 11812 9275 11815
rect 9858 11812 9864 11824
rect 9263 11784 9864 11812
rect 9263 11781 9275 11784
rect 9217 11775 9275 11781
rect 9858 11772 9864 11784
rect 9916 11812 9922 11824
rect 10318 11812 10324 11824
rect 9916 11784 10324 11812
rect 9916 11772 9922 11784
rect 10318 11772 10324 11784
rect 10376 11772 10382 11824
rect 8711 11716 8800 11744
rect 9125 11747 9183 11753
rect 8711 11713 8723 11716
rect 8665 11707 8723 11713
rect 9125 11713 9137 11747
rect 9171 11744 9183 11747
rect 9585 11747 9643 11753
rect 9585 11744 9597 11747
rect 9171 11716 9597 11744
rect 9171 11713 9183 11716
rect 9125 11707 9183 11713
rect 9585 11713 9597 11716
rect 9631 11713 9643 11747
rect 9585 11707 9643 11713
rect 11422 11704 11428 11756
rect 11480 11744 11486 11756
rect 11701 11747 11759 11753
rect 11701 11744 11713 11747
rect 11480 11716 11713 11744
rect 11480 11704 11486 11716
rect 11701 11713 11713 11716
rect 11747 11713 11759 11747
rect 11701 11707 11759 11713
rect 12621 11747 12679 11753
rect 12621 11713 12633 11747
rect 12667 11744 12679 11747
rect 12802 11744 12808 11756
rect 12667 11716 12808 11744
rect 12667 11713 12679 11716
rect 12621 11707 12679 11713
rect 12802 11704 12808 11716
rect 12860 11704 12866 11756
rect 13541 11747 13599 11753
rect 13541 11713 13553 11747
rect 13587 11744 13599 11747
rect 13722 11744 13728 11756
rect 13587 11716 13728 11744
rect 13587 11713 13599 11716
rect 13541 11707 13599 11713
rect 13722 11704 13728 11716
rect 13780 11704 13786 11756
rect 13832 11753 13860 11852
rect 13998 11840 14004 11852
rect 14056 11840 14062 11892
rect 14093 11883 14151 11889
rect 14093 11849 14105 11883
rect 14139 11880 14151 11883
rect 14458 11880 14464 11892
rect 14139 11852 14464 11880
rect 14139 11849 14151 11852
rect 14093 11843 14151 11849
rect 14458 11840 14464 11852
rect 14516 11840 14522 11892
rect 17678 11840 17684 11892
rect 17736 11840 17742 11892
rect 14918 11812 14924 11824
rect 14568 11784 14924 11812
rect 13817 11747 13875 11753
rect 13817 11713 13829 11747
rect 13863 11713 13875 11747
rect 13817 11707 13875 11713
rect 13998 11704 14004 11756
rect 14056 11704 14062 11756
rect 14568 11753 14596 11784
rect 14918 11772 14924 11784
rect 14976 11772 14982 11824
rect 15746 11772 15752 11824
rect 15804 11812 15810 11824
rect 15804 11784 17264 11812
rect 15804 11772 15810 11784
rect 14277 11747 14335 11753
rect 14277 11713 14289 11747
rect 14323 11713 14335 11747
rect 14277 11707 14335 11713
rect 14553 11747 14611 11753
rect 14553 11713 14565 11747
rect 14599 11713 14611 11747
rect 14553 11707 14611 11713
rect 1394 11636 1400 11688
rect 1452 11676 1458 11688
rect 1581 11679 1639 11685
rect 1581 11676 1593 11679
rect 1452 11648 1593 11676
rect 1452 11636 1458 11648
rect 1581 11645 1593 11648
rect 1627 11645 1639 11679
rect 1581 11639 1639 11645
rect 5350 11636 5356 11688
rect 5408 11676 5414 11688
rect 5629 11679 5687 11685
rect 5629 11676 5641 11679
rect 5408 11648 5641 11676
rect 5408 11636 5414 11648
rect 5629 11645 5641 11648
rect 5675 11645 5687 11679
rect 5629 11639 5687 11645
rect 9309 11679 9367 11685
rect 9309 11645 9321 11679
rect 9355 11645 9367 11679
rect 9309 11639 9367 11645
rect 4614 11568 4620 11620
rect 4672 11608 4678 11620
rect 5077 11611 5135 11617
rect 5077 11608 5089 11611
rect 4672 11580 5089 11608
rect 4672 11568 4678 11580
rect 5077 11577 5089 11580
rect 5123 11577 5135 11611
rect 5077 11571 5135 11577
rect 5902 11568 5908 11620
rect 5960 11608 5966 11620
rect 6822 11608 6828 11620
rect 5960 11580 6828 11608
rect 5960 11568 5966 11580
rect 6822 11568 6828 11580
rect 6880 11568 6886 11620
rect 8662 11568 8668 11620
rect 8720 11608 8726 11620
rect 9324 11608 9352 11639
rect 9398 11636 9404 11688
rect 9456 11676 9462 11688
rect 10137 11679 10195 11685
rect 10137 11676 10149 11679
rect 9456 11648 10149 11676
rect 9456 11636 9462 11648
rect 10137 11645 10149 11648
rect 10183 11645 10195 11679
rect 14292 11676 14320 11707
rect 14642 11704 14648 11756
rect 14700 11744 14706 11756
rect 14737 11747 14795 11753
rect 14737 11744 14749 11747
rect 14700 11716 14749 11744
rect 14700 11704 14706 11716
rect 14737 11713 14749 11716
rect 14783 11744 14795 11747
rect 15010 11744 15016 11756
rect 14783 11716 15016 11744
rect 14783 11713 14795 11716
rect 14737 11707 14795 11713
rect 15010 11704 15016 11716
rect 15068 11704 15074 11756
rect 15565 11747 15623 11753
rect 15565 11713 15577 11747
rect 15611 11713 15623 11747
rect 15565 11707 15623 11713
rect 16485 11747 16543 11753
rect 16485 11713 16497 11747
rect 16531 11744 16543 11747
rect 17037 11747 17095 11753
rect 17037 11744 17049 11747
rect 16531 11716 17049 11744
rect 16531 11713 16543 11716
rect 16485 11707 16543 11713
rect 17037 11713 17049 11716
rect 17083 11713 17095 11747
rect 17037 11707 17095 11713
rect 10137 11639 10195 11645
rect 13740 11648 14320 11676
rect 13740 11620 13768 11648
rect 8720 11580 9352 11608
rect 8720 11568 8726 11580
rect 2866 11500 2872 11552
rect 2924 11540 2930 11552
rect 2961 11543 3019 11549
rect 2961 11540 2973 11543
rect 2924 11512 2973 11540
rect 2924 11500 2930 11512
rect 2961 11509 2973 11512
rect 3007 11509 3019 11543
rect 2961 11503 3019 11509
rect 4985 11543 5043 11549
rect 4985 11509 4997 11543
rect 5031 11540 5043 11543
rect 5350 11540 5356 11552
rect 5031 11512 5356 11540
rect 5031 11509 5043 11512
rect 4985 11503 5043 11509
rect 5350 11500 5356 11512
rect 5408 11500 5414 11552
rect 6362 11500 6368 11552
rect 6420 11500 6426 11552
rect 8478 11500 8484 11552
rect 8536 11500 8542 11552
rect 9324 11540 9352 11580
rect 13078 11568 13084 11620
rect 13136 11568 13142 11620
rect 13722 11568 13728 11620
rect 13780 11568 13786 11620
rect 15580 11608 15608 11707
rect 17236 11688 17264 11784
rect 17494 11704 17500 11756
rect 17552 11704 17558 11756
rect 15933 11679 15991 11685
rect 15933 11645 15945 11679
rect 15979 11676 15991 11679
rect 16206 11676 16212 11688
rect 15979 11648 16212 11676
rect 15979 11645 15991 11648
rect 15933 11639 15991 11645
rect 16206 11636 16212 11648
rect 16264 11636 16270 11688
rect 17126 11636 17132 11688
rect 17184 11636 17190 11688
rect 17218 11636 17224 11688
rect 17276 11636 17282 11688
rect 16669 11611 16727 11617
rect 16669 11608 16681 11611
rect 15580 11580 16681 11608
rect 16669 11577 16681 11580
rect 16715 11577 16727 11611
rect 16669 11571 16727 11577
rect 11146 11540 11152 11552
rect 9324 11512 11152 11540
rect 11146 11500 11152 11512
rect 11204 11500 11210 11552
rect 11517 11543 11575 11549
rect 11517 11509 11529 11543
rect 11563 11540 11575 11543
rect 12250 11540 12256 11552
rect 11563 11512 12256 11540
rect 11563 11509 11575 11512
rect 11517 11503 11575 11509
rect 12250 11500 12256 11512
rect 12308 11500 12314 11552
rect 12618 11500 12624 11552
rect 12676 11540 12682 11552
rect 12713 11543 12771 11549
rect 12713 11540 12725 11543
rect 12676 11512 12725 11540
rect 12676 11500 12682 11512
rect 12713 11509 12725 11512
rect 12759 11509 12771 11543
rect 12713 11503 12771 11509
rect 13357 11543 13415 11549
rect 13357 11509 13369 11543
rect 13403 11540 13415 11543
rect 13538 11540 13544 11552
rect 13403 11512 13544 11540
rect 13403 11509 13415 11512
rect 13357 11503 13415 11509
rect 13538 11500 13544 11512
rect 13596 11500 13602 11552
rect 15746 11500 15752 11552
rect 15804 11500 15810 11552
rect 1104 11450 18124 11472
rect 1104 11398 3077 11450
rect 3129 11398 3141 11450
rect 3193 11398 3205 11450
rect 3257 11398 3269 11450
rect 3321 11398 3333 11450
rect 3385 11398 7332 11450
rect 7384 11398 7396 11450
rect 7448 11398 7460 11450
rect 7512 11398 7524 11450
rect 7576 11398 7588 11450
rect 7640 11398 11587 11450
rect 11639 11398 11651 11450
rect 11703 11398 11715 11450
rect 11767 11398 11779 11450
rect 11831 11398 11843 11450
rect 11895 11398 15842 11450
rect 15894 11398 15906 11450
rect 15958 11398 15970 11450
rect 16022 11398 16034 11450
rect 16086 11398 16098 11450
rect 16150 11398 18124 11450
rect 1104 11376 18124 11398
rect 2038 11296 2044 11348
rect 2096 11296 2102 11348
rect 3878 11296 3884 11348
rect 3936 11336 3942 11348
rect 3973 11339 4031 11345
rect 3973 11336 3985 11339
rect 3936 11308 3985 11336
rect 3936 11296 3942 11308
rect 3973 11305 3985 11308
rect 4019 11305 4031 11339
rect 3973 11299 4031 11305
rect 5350 11296 5356 11348
rect 5408 11296 5414 11348
rect 6546 11296 6552 11348
rect 6604 11336 6610 11348
rect 9766 11336 9772 11348
rect 6604 11308 9772 11336
rect 6604 11296 6610 11308
rect 4249 11271 4307 11277
rect 4249 11237 4261 11271
rect 4295 11237 4307 11271
rect 4249 11231 4307 11237
rect 2314 11160 2320 11212
rect 2372 11200 2378 11212
rect 2593 11203 2651 11209
rect 2593 11200 2605 11203
rect 2372 11172 2605 11200
rect 2372 11160 2378 11172
rect 2593 11169 2605 11172
rect 2639 11169 2651 11203
rect 2593 11163 2651 11169
rect 1946 11092 1952 11144
rect 2004 11092 2010 11144
rect 2406 11092 2412 11144
rect 2464 11092 2470 11144
rect 2608 11132 2636 11163
rect 2958 11160 2964 11212
rect 3016 11160 3022 11212
rect 3050 11132 3056 11144
rect 2608 11104 3056 11132
rect 3050 11092 3056 11104
rect 3108 11092 3114 11144
rect 4157 11135 4215 11141
rect 4157 11101 4169 11135
rect 4203 11132 4215 11135
rect 4264 11132 4292 11231
rect 5534 11228 5540 11280
rect 5592 11268 5598 11280
rect 6086 11268 6092 11280
rect 5592 11240 6092 11268
rect 5592 11228 5598 11240
rect 6086 11228 6092 11240
rect 6144 11228 6150 11280
rect 4798 11160 4804 11212
rect 4856 11160 4862 11212
rect 5000 11172 6592 11200
rect 4203 11104 4292 11132
rect 4203 11101 4215 11104
rect 4157 11095 4215 11101
rect 4614 11092 4620 11144
rect 4672 11092 4678 11144
rect 4706 11092 4712 11144
rect 4764 11132 4770 11144
rect 5000 11132 5028 11172
rect 4764 11104 5028 11132
rect 4764 11092 4770 11104
rect 5074 11092 5080 11144
rect 5132 11092 5138 11144
rect 5534 11092 5540 11144
rect 5592 11132 5598 11144
rect 5810 11141 5816 11144
rect 5629 11135 5687 11141
rect 5629 11132 5641 11135
rect 5592 11104 5641 11132
rect 5592 11092 5598 11104
rect 5629 11101 5641 11104
rect 5675 11101 5687 11135
rect 5629 11095 5687 11101
rect 5777 11135 5816 11141
rect 5777 11101 5789 11135
rect 5777 11095 5816 11101
rect 5810 11092 5816 11095
rect 5868 11092 5874 11144
rect 6135 11135 6193 11141
rect 6135 11101 6147 11135
rect 6181 11132 6193 11135
rect 6457 11135 6515 11141
rect 6457 11132 6469 11135
rect 6181 11104 6469 11132
rect 6181 11101 6193 11104
rect 6135 11095 6193 11101
rect 6457 11101 6469 11104
rect 6503 11101 6515 11135
rect 6457 11095 6515 11101
rect 1486 11024 1492 11076
rect 1544 11024 1550 11076
rect 1673 11067 1731 11073
rect 1673 11033 1685 11067
rect 1719 11064 1731 11067
rect 1719 11036 2544 11064
rect 1719 11033 1731 11036
rect 1673 11027 1731 11033
rect 1762 10956 1768 11008
rect 1820 10956 1826 11008
rect 2516 11005 2544 11036
rect 2866 11024 2872 11076
rect 2924 11064 2930 11076
rect 5905 11067 5963 11073
rect 5905 11064 5917 11067
rect 2924 11036 3280 11064
rect 2924 11024 2930 11036
rect 3252 11008 3280 11036
rect 3620 11036 5917 11064
rect 2501 10999 2559 11005
rect 2501 10965 2513 10999
rect 2547 10996 2559 10999
rect 2682 10996 2688 11008
rect 2547 10968 2688 10996
rect 2547 10965 2559 10968
rect 2501 10959 2559 10965
rect 2682 10956 2688 10968
rect 2740 10956 2746 11008
rect 3142 10956 3148 11008
rect 3200 10956 3206 11008
rect 3234 10956 3240 11008
rect 3292 10956 3298 11008
rect 3620 11005 3648 11036
rect 5905 11033 5917 11036
rect 5951 11033 5963 11067
rect 5905 11027 5963 11033
rect 5994 11024 6000 11076
rect 6052 11024 6058 11076
rect 6564 11064 6592 11172
rect 6656 11141 6684 11308
rect 9766 11296 9772 11308
rect 9824 11296 9830 11348
rect 13078 11296 13084 11348
rect 13136 11336 13142 11348
rect 14090 11336 14096 11348
rect 13136 11308 14096 11336
rect 13136 11296 13142 11308
rect 14090 11296 14096 11308
rect 14148 11296 14154 11348
rect 12802 11228 12808 11280
rect 12860 11268 12866 11280
rect 14366 11268 14372 11280
rect 12860 11240 14372 11268
rect 12860 11228 12866 11240
rect 14366 11228 14372 11240
rect 14424 11228 14430 11280
rect 14918 11228 14924 11280
rect 14976 11268 14982 11280
rect 14976 11240 16160 11268
rect 14976 11228 14982 11240
rect 7024 11172 7696 11200
rect 7024 11144 7052 11172
rect 6641 11135 6699 11141
rect 6641 11101 6653 11135
rect 6687 11101 6699 11135
rect 6641 11095 6699 11101
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11132 6975 11135
rect 7006 11132 7012 11144
rect 6963 11104 7012 11132
rect 6963 11101 6975 11104
rect 6917 11095 6975 11101
rect 7006 11092 7012 11104
rect 7064 11092 7070 11144
rect 7101 11135 7159 11141
rect 7101 11101 7113 11135
rect 7147 11132 7159 11135
rect 7190 11132 7196 11144
rect 7147 11104 7196 11132
rect 7147 11101 7159 11104
rect 7101 11095 7159 11101
rect 7190 11092 7196 11104
rect 7248 11092 7254 11144
rect 7668 11132 7696 11172
rect 7834 11160 7840 11212
rect 7892 11160 7898 11212
rect 15010 11160 15016 11212
rect 15068 11200 15074 11212
rect 16132 11209 16160 11240
rect 16206 11228 16212 11280
rect 16264 11268 16270 11280
rect 16393 11271 16451 11277
rect 16393 11268 16405 11271
rect 16264 11240 16405 11268
rect 16264 11228 16270 11240
rect 16393 11237 16405 11240
rect 16439 11237 16451 11271
rect 16393 11231 16451 11237
rect 15289 11203 15347 11209
rect 15289 11200 15301 11203
rect 15068 11172 15301 11200
rect 15068 11160 15074 11172
rect 15289 11169 15301 11172
rect 15335 11169 15347 11203
rect 15289 11163 15347 11169
rect 16117 11203 16175 11209
rect 16117 11169 16129 11203
rect 16163 11169 16175 11203
rect 16117 11163 16175 11169
rect 8665 11135 8723 11141
rect 8665 11132 8677 11135
rect 7668 11104 8677 11132
rect 8665 11101 8677 11104
rect 8711 11101 8723 11135
rect 8665 11095 8723 11101
rect 9493 11135 9551 11141
rect 9493 11101 9505 11135
rect 9539 11132 9551 11135
rect 9674 11132 9680 11144
rect 9539 11104 9680 11132
rect 9539 11101 9551 11104
rect 9493 11095 9551 11101
rect 9674 11092 9680 11104
rect 9732 11092 9738 11144
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11132 9827 11135
rect 11241 11135 11299 11141
rect 11241 11132 11253 11135
rect 9815 11104 11253 11132
rect 9815 11101 9827 11104
rect 9769 11095 9827 11101
rect 11241 11101 11253 11104
rect 11287 11132 11299 11135
rect 11330 11132 11336 11144
rect 11287 11104 11336 11132
rect 11287 11101 11299 11104
rect 11241 11095 11299 11101
rect 11330 11092 11336 11104
rect 11388 11092 11394 11144
rect 11508 11135 11566 11141
rect 11508 11101 11520 11135
rect 11554 11132 11566 11135
rect 12250 11132 12256 11144
rect 11554 11104 12256 11132
rect 11554 11101 11566 11104
rect 11508 11095 11566 11101
rect 12250 11092 12256 11104
rect 12308 11092 12314 11144
rect 12618 11092 12624 11144
rect 12676 11132 12682 11144
rect 13265 11135 13323 11141
rect 13265 11132 13277 11135
rect 12676 11104 13277 11132
rect 12676 11092 12682 11104
rect 13265 11101 13277 11104
rect 13311 11101 13323 11135
rect 13265 11095 13323 11101
rect 15105 11135 15163 11141
rect 15105 11101 15117 11135
rect 15151 11132 15163 11135
rect 15933 11135 15991 11141
rect 15933 11132 15945 11135
rect 15151 11104 15945 11132
rect 15151 11101 15163 11104
rect 15105 11095 15163 11101
rect 15933 11101 15945 11104
rect 15979 11132 15991 11135
rect 16224 11132 16252 11228
rect 15979 11104 16252 11132
rect 15979 11101 15991 11104
rect 15933 11095 15991 11101
rect 16390 11092 16396 11144
rect 16448 11132 16454 11144
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 16448 11104 17785 11132
rect 16448 11092 16454 11104
rect 17773 11101 17785 11104
rect 17819 11101 17831 11135
rect 17773 11095 17831 11101
rect 7653 11067 7711 11073
rect 7653 11064 7665 11067
rect 6564 11036 7665 11064
rect 7116 11008 7144 11036
rect 7653 11033 7665 11036
rect 7699 11033 7711 11067
rect 7653 11027 7711 11033
rect 7745 11067 7803 11073
rect 7745 11033 7757 11067
rect 7791 11064 7803 11067
rect 8113 11067 8171 11073
rect 8113 11064 8125 11067
rect 7791 11036 8125 11064
rect 7791 11033 7803 11036
rect 7745 11027 7803 11033
rect 8113 11033 8125 11036
rect 8159 11033 8171 11067
rect 10014 11067 10072 11073
rect 10014 11064 10026 11067
rect 8113 11027 8171 11033
rect 9692 11036 10026 11064
rect 3605 10999 3663 11005
rect 3605 10965 3617 10999
rect 3651 10965 3663 10999
rect 3605 10959 3663 10965
rect 5534 10956 5540 11008
rect 5592 10956 5598 11008
rect 6270 10956 6276 11008
rect 6328 10956 6334 11008
rect 7098 10956 7104 11008
rect 7156 10956 7162 11008
rect 7190 10956 7196 11008
rect 7248 10996 7254 11008
rect 9692 11005 9720 11036
rect 10014 11033 10026 11036
rect 10060 11033 10072 11067
rect 10014 11027 10072 11033
rect 12066 11024 12072 11076
rect 12124 11064 12130 11076
rect 12713 11067 12771 11073
rect 12713 11064 12725 11067
rect 12124 11036 12725 11064
rect 12124 11024 12130 11036
rect 12713 11033 12725 11036
rect 12759 11033 12771 11067
rect 12713 11027 12771 11033
rect 15197 11067 15255 11073
rect 15197 11033 15209 11067
rect 15243 11064 15255 11067
rect 15243 11036 15700 11064
rect 15243 11033 15255 11036
rect 15197 11027 15255 11033
rect 7285 10999 7343 11005
rect 7285 10996 7297 10999
rect 7248 10968 7297 10996
rect 7248 10956 7254 10968
rect 7285 10965 7297 10968
rect 7331 10965 7343 10999
rect 7285 10959 7343 10965
rect 9677 10999 9735 11005
rect 9677 10965 9689 10999
rect 9723 10965 9735 10999
rect 9677 10959 9735 10965
rect 11149 10999 11207 11005
rect 11149 10965 11161 10999
rect 11195 10996 11207 10999
rect 11330 10996 11336 11008
rect 11195 10968 11336 10996
rect 11195 10965 11207 10968
rect 11149 10959 11207 10965
rect 11330 10956 11336 10968
rect 11388 10956 11394 11008
rect 12618 10956 12624 11008
rect 12676 10956 12682 11008
rect 14182 10956 14188 11008
rect 14240 10996 14246 11008
rect 14737 10999 14795 11005
rect 14737 10996 14749 10999
rect 14240 10968 14749 10996
rect 14240 10956 14246 10968
rect 14737 10965 14749 10968
rect 14783 10965 14795 10999
rect 14737 10959 14795 10965
rect 15102 10956 15108 11008
rect 15160 10996 15166 11008
rect 15212 10996 15240 11027
rect 15160 10968 15240 10996
rect 15160 10956 15166 10968
rect 15562 10956 15568 11008
rect 15620 10956 15626 11008
rect 15672 10996 15700 11036
rect 15746 11024 15752 11076
rect 15804 11064 15810 11076
rect 17506 11067 17564 11073
rect 17506 11064 17518 11067
rect 15804 11036 17518 11064
rect 15804 11024 15810 11036
rect 17506 11033 17518 11036
rect 17552 11033 17564 11067
rect 17506 11027 17564 11033
rect 16025 10999 16083 11005
rect 16025 10996 16037 10999
rect 15672 10968 16037 10996
rect 16025 10965 16037 10968
rect 16071 10996 16083 10999
rect 16850 10996 16856 11008
rect 16071 10968 16856 10996
rect 16071 10965 16083 10968
rect 16025 10959 16083 10965
rect 16850 10956 16856 10968
rect 16908 10956 16914 11008
rect 1104 10906 18124 10928
rect 1104 10854 3737 10906
rect 3789 10854 3801 10906
rect 3853 10854 3865 10906
rect 3917 10854 3929 10906
rect 3981 10854 3993 10906
rect 4045 10854 7992 10906
rect 8044 10854 8056 10906
rect 8108 10854 8120 10906
rect 8172 10854 8184 10906
rect 8236 10854 8248 10906
rect 8300 10854 12247 10906
rect 12299 10854 12311 10906
rect 12363 10854 12375 10906
rect 12427 10854 12439 10906
rect 12491 10854 12503 10906
rect 12555 10854 16502 10906
rect 16554 10854 16566 10906
rect 16618 10854 16630 10906
rect 16682 10854 16694 10906
rect 16746 10854 16758 10906
rect 16810 10854 18124 10906
rect 1104 10832 18124 10854
rect 2777 10795 2835 10801
rect 2777 10761 2789 10795
rect 2823 10792 2835 10795
rect 3142 10792 3148 10804
rect 2823 10764 3148 10792
rect 2823 10761 2835 10764
rect 2777 10755 2835 10761
rect 3142 10752 3148 10764
rect 3200 10752 3206 10804
rect 3234 10752 3240 10804
rect 3292 10792 3298 10804
rect 3697 10795 3755 10801
rect 3697 10792 3709 10795
rect 3292 10764 3709 10792
rect 3292 10752 3298 10764
rect 3697 10761 3709 10764
rect 3743 10761 3755 10795
rect 3697 10755 3755 10761
rect 4065 10795 4123 10801
rect 4065 10761 4077 10795
rect 4111 10761 4123 10795
rect 4065 10755 4123 10761
rect 1664 10727 1722 10733
rect 1664 10693 1676 10727
rect 1710 10724 1722 10727
rect 1762 10724 1768 10736
rect 1710 10696 1768 10724
rect 1710 10693 1722 10696
rect 1664 10687 1722 10693
rect 1762 10684 1768 10696
rect 1820 10684 1826 10736
rect 4080 10724 4108 10755
rect 5534 10752 5540 10804
rect 5592 10792 5598 10804
rect 5592 10764 5948 10792
rect 5592 10752 5598 10764
rect 5920 10733 5948 10764
rect 7006 10752 7012 10804
rect 7064 10792 7070 10804
rect 7929 10795 7987 10801
rect 7929 10792 7941 10795
rect 7064 10764 7941 10792
rect 7064 10752 7070 10764
rect 7929 10761 7941 10764
rect 7975 10761 7987 10795
rect 7929 10755 7987 10761
rect 9398 10752 9404 10804
rect 9456 10752 9462 10804
rect 10778 10752 10784 10804
rect 10836 10752 10842 10804
rect 11422 10752 11428 10804
rect 11480 10792 11486 10804
rect 11701 10795 11759 10801
rect 11701 10792 11713 10795
rect 11480 10764 11713 10792
rect 11480 10752 11486 10764
rect 11701 10761 11713 10764
rect 11747 10761 11759 10795
rect 11701 10755 11759 10761
rect 12066 10752 12072 10804
rect 12124 10752 12130 10804
rect 13262 10752 13268 10804
rect 13320 10752 13326 10804
rect 13446 10752 13452 10804
rect 13504 10792 13510 10804
rect 13725 10795 13783 10801
rect 13725 10792 13737 10795
rect 13504 10764 13737 10792
rect 13504 10752 13510 10764
rect 13725 10761 13737 10764
rect 13771 10761 13783 10795
rect 13725 10755 13783 10761
rect 13817 10795 13875 10801
rect 13817 10761 13829 10795
rect 13863 10792 13875 10795
rect 13906 10792 13912 10804
rect 13863 10764 13912 10792
rect 13863 10761 13875 10764
rect 13817 10755 13875 10761
rect 13906 10752 13912 10764
rect 13964 10752 13970 10804
rect 15562 10792 15568 10804
rect 14016 10764 15568 10792
rect 5813 10727 5871 10733
rect 5813 10724 5825 10727
rect 4080 10696 5825 10724
rect 5813 10693 5825 10696
rect 5859 10693 5871 10727
rect 5813 10687 5871 10693
rect 5905 10727 5963 10733
rect 5905 10693 5917 10727
rect 5951 10693 5963 10727
rect 6914 10724 6920 10736
rect 5905 10687 5963 10693
rect 6564 10696 6920 10724
rect 1394 10616 1400 10668
rect 1452 10616 1458 10668
rect 3142 10616 3148 10668
rect 3200 10656 3206 10668
rect 3605 10659 3663 10665
rect 3605 10656 3617 10659
rect 3200 10628 3617 10656
rect 3200 10616 3206 10628
rect 3605 10625 3617 10628
rect 3651 10656 3663 10659
rect 4709 10659 4767 10665
rect 4709 10656 4721 10659
rect 3651 10628 4721 10656
rect 3651 10625 3663 10628
rect 3605 10619 3663 10625
rect 4709 10625 4721 10628
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 4985 10659 5043 10665
rect 4985 10625 4997 10659
rect 5031 10656 5043 10659
rect 5258 10656 5264 10668
rect 5031 10628 5264 10656
rect 5031 10625 5043 10628
rect 4985 10619 5043 10625
rect 5258 10616 5264 10628
rect 5316 10616 5322 10668
rect 5534 10616 5540 10668
rect 5592 10616 5598 10668
rect 5718 10665 5724 10668
rect 5685 10659 5724 10665
rect 5685 10625 5697 10659
rect 5685 10619 5724 10625
rect 5718 10616 5724 10619
rect 5776 10616 5782 10668
rect 6043 10659 6101 10665
rect 6043 10625 6055 10659
rect 6089 10656 6101 10659
rect 6362 10656 6368 10668
rect 6089 10628 6368 10656
rect 6089 10625 6101 10628
rect 6043 10619 6101 10625
rect 6362 10616 6368 10628
rect 6420 10616 6426 10668
rect 6564 10665 6592 10696
rect 6914 10684 6920 10696
rect 6972 10724 6978 10736
rect 8288 10727 8346 10733
rect 6972 10696 8064 10724
rect 6972 10684 6978 10696
rect 6822 10665 6828 10668
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10625 6607 10659
rect 6549 10619 6607 10625
rect 6816 10619 6828 10665
rect 6822 10616 6828 10619
rect 6880 10616 6886 10668
rect 8036 10665 8064 10696
rect 8288 10693 8300 10727
rect 8334 10724 8346 10727
rect 8478 10724 8484 10736
rect 8334 10696 8484 10724
rect 8334 10693 8346 10696
rect 8288 10687 8346 10693
rect 8478 10684 8484 10696
rect 8536 10684 8542 10736
rect 10962 10684 10968 10736
rect 11020 10724 11026 10736
rect 12161 10727 12219 10733
rect 12161 10724 12173 10727
rect 11020 10696 12173 10724
rect 11020 10684 11026 10696
rect 12161 10693 12173 10696
rect 12207 10724 12219 10727
rect 13280 10724 13308 10752
rect 12207 10696 12940 10724
rect 12207 10693 12219 10696
rect 12161 10687 12219 10693
rect 8021 10659 8079 10665
rect 8021 10625 8033 10659
rect 8067 10625 8079 10659
rect 8021 10619 8079 10625
rect 9490 10616 9496 10668
rect 9548 10616 9554 10668
rect 11146 10616 11152 10668
rect 11204 10656 11210 10668
rect 11974 10656 11980 10668
rect 11204 10628 11980 10656
rect 11204 10616 11210 10628
rect 11974 10616 11980 10628
rect 12032 10656 12038 10668
rect 12529 10659 12587 10665
rect 12032 10628 12296 10656
rect 12032 10616 12038 10628
rect 12268 10600 12296 10628
rect 12529 10625 12541 10659
rect 12575 10656 12587 10659
rect 12710 10656 12716 10668
rect 12575 10628 12716 10656
rect 12575 10625 12587 10628
rect 12529 10619 12587 10625
rect 12710 10616 12716 10628
rect 12768 10616 12774 10668
rect 2774 10548 2780 10600
rect 2832 10588 2838 10600
rect 3418 10588 3424 10600
rect 2832 10560 3424 10588
rect 2832 10548 2838 10560
rect 3418 10548 3424 10560
rect 3476 10548 3482 10600
rect 12250 10548 12256 10600
rect 12308 10548 12314 10600
rect 5445 10523 5503 10529
rect 5445 10489 5457 10523
rect 5491 10520 5503 10523
rect 5994 10520 6000 10532
rect 5491 10492 6000 10520
rect 5491 10489 5503 10492
rect 5445 10483 5503 10489
rect 5994 10480 6000 10492
rect 6052 10480 6058 10532
rect 12912 10520 12940 10696
rect 13096 10696 13308 10724
rect 13357 10727 13415 10733
rect 13096 10668 13124 10696
rect 13357 10693 13369 10727
rect 13403 10724 13415 10727
rect 14016 10724 14044 10764
rect 15562 10752 15568 10764
rect 15620 10752 15626 10804
rect 13403 10696 14044 10724
rect 13403 10693 13415 10696
rect 13357 10687 13415 10693
rect 14090 10684 14096 10736
rect 14148 10684 14154 10736
rect 14182 10684 14188 10736
rect 14240 10684 14246 10736
rect 13078 10616 13084 10668
rect 13136 10616 13142 10668
rect 13262 10665 13268 10668
rect 13229 10659 13268 10665
rect 13229 10625 13241 10659
rect 13229 10619 13268 10625
rect 13262 10616 13268 10619
rect 13320 10616 13326 10668
rect 13449 10659 13507 10665
rect 13449 10625 13461 10659
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 12989 10591 13047 10597
rect 12989 10557 13001 10591
rect 13035 10588 13047 10591
rect 13464 10588 13492 10619
rect 13538 10616 13544 10668
rect 13596 10665 13602 10668
rect 13596 10656 13604 10665
rect 13596 10628 13641 10656
rect 13596 10619 13604 10628
rect 13596 10616 13602 10619
rect 13906 10616 13912 10668
rect 13964 10665 13970 10668
rect 13964 10659 14013 10665
rect 13964 10625 13967 10659
rect 14001 10625 14013 10659
rect 13964 10619 14013 10625
rect 13964 10616 13970 10619
rect 14274 10616 14280 10668
rect 14332 10665 14338 10668
rect 14332 10659 14371 10665
rect 14359 10625 14371 10659
rect 14332 10619 14371 10625
rect 14461 10659 14519 10665
rect 14461 10625 14473 10659
rect 14507 10656 14519 10659
rect 14550 10656 14556 10668
rect 14507 10628 14556 10656
rect 14507 10625 14519 10628
rect 14461 10619 14519 10625
rect 14332 10616 14338 10619
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 14737 10659 14795 10665
rect 14737 10625 14749 10659
rect 14783 10656 14795 10659
rect 14826 10656 14832 10668
rect 14783 10628 14832 10656
rect 14783 10625 14795 10628
rect 14737 10619 14795 10625
rect 14826 10616 14832 10628
rect 14884 10616 14890 10668
rect 16206 10616 16212 10668
rect 16264 10665 16270 10668
rect 16264 10619 16276 10665
rect 16264 10616 16270 10619
rect 16390 10616 16396 10668
rect 16448 10656 16454 10668
rect 16485 10659 16543 10665
rect 16485 10656 16497 10659
rect 16448 10628 16497 10656
rect 16448 10616 16454 10628
rect 16485 10625 16497 10628
rect 16531 10625 16543 10659
rect 16485 10619 16543 10625
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10656 17095 10659
rect 17494 10656 17500 10668
rect 17083 10628 17500 10656
rect 17083 10625 17095 10628
rect 17037 10619 17095 10625
rect 17494 10616 17500 10628
rect 17552 10616 17558 10668
rect 17678 10616 17684 10668
rect 17736 10616 17742 10668
rect 17126 10588 17132 10600
rect 13035 10560 13492 10588
rect 16500 10560 17132 10588
rect 13035 10557 13047 10560
rect 12989 10551 13047 10557
rect 14458 10520 14464 10532
rect 12912 10492 14464 10520
rect 14458 10480 14464 10492
rect 14516 10520 14522 10532
rect 14516 10492 15056 10520
rect 14516 10480 14522 10492
rect 4154 10412 4160 10464
rect 4212 10412 4218 10464
rect 5261 10455 5319 10461
rect 5261 10421 5273 10455
rect 5307 10452 5319 10455
rect 5350 10452 5356 10464
rect 5307 10424 5356 10452
rect 5307 10421 5319 10424
rect 5261 10415 5319 10421
rect 5350 10412 5356 10424
rect 5408 10412 5414 10464
rect 6181 10455 6239 10461
rect 6181 10421 6193 10455
rect 6227 10452 6239 10455
rect 7834 10452 7840 10464
rect 6227 10424 7840 10452
rect 6227 10421 6239 10424
rect 6181 10415 6239 10421
rect 7834 10412 7840 10424
rect 7892 10412 7898 10464
rect 12618 10412 12624 10464
rect 12676 10412 12682 10464
rect 14550 10412 14556 10464
rect 14608 10412 14614 10464
rect 15028 10452 15056 10492
rect 15102 10480 15108 10532
rect 15160 10480 15166 10532
rect 16500 10452 16528 10560
rect 17126 10548 17132 10560
rect 17184 10548 17190 10600
rect 17310 10548 17316 10600
rect 17368 10548 17374 10600
rect 17144 10520 17172 10548
rect 17497 10523 17555 10529
rect 17497 10520 17509 10523
rect 17144 10492 17509 10520
rect 17497 10489 17509 10492
rect 17543 10489 17555 10523
rect 17497 10483 17555 10489
rect 15028 10424 16528 10452
rect 16666 10412 16672 10464
rect 16724 10412 16730 10464
rect 1104 10362 18124 10384
rect 1104 10310 3077 10362
rect 3129 10310 3141 10362
rect 3193 10310 3205 10362
rect 3257 10310 3269 10362
rect 3321 10310 3333 10362
rect 3385 10310 7332 10362
rect 7384 10310 7396 10362
rect 7448 10310 7460 10362
rect 7512 10310 7524 10362
rect 7576 10310 7588 10362
rect 7640 10310 11587 10362
rect 11639 10310 11651 10362
rect 11703 10310 11715 10362
rect 11767 10310 11779 10362
rect 11831 10310 11843 10362
rect 11895 10310 15842 10362
rect 15894 10310 15906 10362
rect 15958 10310 15970 10362
rect 16022 10310 16034 10362
rect 16086 10310 16098 10362
rect 16150 10310 18124 10362
rect 1104 10288 18124 10310
rect 1210 10208 1216 10260
rect 1268 10248 1274 10260
rect 1489 10251 1547 10257
rect 1489 10248 1501 10251
rect 1268 10220 1501 10248
rect 1268 10208 1274 10220
rect 1489 10217 1501 10220
rect 1535 10217 1547 10251
rect 1489 10211 1547 10217
rect 1946 10208 1952 10260
rect 2004 10248 2010 10260
rect 2225 10251 2283 10257
rect 2225 10248 2237 10251
rect 2004 10220 2237 10248
rect 2004 10208 2010 10220
rect 2225 10217 2237 10220
rect 2271 10217 2283 10251
rect 2225 10211 2283 10217
rect 6822 10208 6828 10260
rect 6880 10248 6886 10260
rect 7285 10251 7343 10257
rect 7285 10248 7297 10251
rect 6880 10220 7297 10248
rect 6880 10208 6886 10220
rect 7285 10217 7297 10220
rect 7331 10217 7343 10251
rect 7285 10211 7343 10217
rect 9674 10208 9680 10260
rect 9732 10248 9738 10260
rect 9953 10251 10011 10257
rect 9953 10248 9965 10251
rect 9732 10220 9965 10248
rect 9732 10208 9738 10220
rect 9953 10217 9965 10220
rect 9999 10217 10011 10251
rect 12253 10251 12311 10257
rect 12253 10248 12265 10251
rect 9953 10211 10011 10217
rect 10520 10220 12265 10248
rect 2590 10140 2596 10192
rect 2648 10140 2654 10192
rect 9766 10140 9772 10192
rect 9824 10180 9830 10192
rect 10520 10180 10548 10220
rect 12253 10217 12265 10220
rect 12299 10248 12311 10251
rect 12618 10248 12624 10260
rect 12299 10220 12624 10248
rect 12299 10217 12311 10220
rect 12253 10211 12311 10217
rect 12618 10208 12624 10220
rect 12676 10208 12682 10260
rect 12802 10208 12808 10260
rect 12860 10208 12866 10260
rect 13906 10208 13912 10260
rect 13964 10208 13970 10260
rect 14826 10208 14832 10260
rect 14884 10208 14890 10260
rect 16025 10251 16083 10257
rect 16025 10217 16037 10251
rect 16071 10248 16083 10251
rect 16206 10248 16212 10260
rect 16071 10220 16212 10248
rect 16071 10217 16083 10220
rect 16025 10211 16083 10217
rect 16206 10208 16212 10220
rect 16264 10208 16270 10260
rect 17494 10208 17500 10260
rect 17552 10208 17558 10260
rect 9824 10152 10548 10180
rect 10612 10152 14320 10180
rect 9824 10140 9830 10152
rect 2608 10112 2636 10140
rect 2777 10115 2835 10121
rect 2777 10112 2789 10115
rect 2608 10084 2789 10112
rect 2777 10081 2789 10084
rect 2823 10081 2835 10115
rect 2777 10075 2835 10081
rect 7926 10072 7932 10124
rect 7984 10112 7990 10124
rect 8386 10112 8392 10124
rect 7984 10084 8392 10112
rect 7984 10072 7990 10084
rect 8386 10072 8392 10084
rect 8444 10112 8450 10124
rect 10612 10121 10640 10152
rect 10597 10115 10655 10121
rect 10597 10112 10609 10115
rect 8444 10084 10609 10112
rect 8444 10072 8450 10084
rect 10597 10081 10609 10084
rect 10643 10081 10655 10115
rect 10597 10075 10655 10081
rect 11330 10072 11336 10124
rect 11388 10072 11394 10124
rect 14292 10121 14320 10152
rect 14277 10115 14335 10121
rect 12268 10084 13768 10112
rect 1673 10047 1731 10053
rect 1673 10013 1685 10047
rect 1719 10013 1731 10047
rect 1673 10007 1731 10013
rect 1688 9976 1716 10007
rect 2038 10004 2044 10056
rect 2096 10004 2102 10056
rect 2593 10047 2651 10053
rect 2593 10013 2605 10047
rect 2639 10044 2651 10047
rect 4154 10044 4160 10056
rect 2639 10016 4160 10044
rect 2639 10013 2651 10016
rect 2593 10007 2651 10013
rect 4154 10004 4160 10016
rect 4212 10004 4218 10056
rect 7190 10004 7196 10056
rect 7248 10044 7254 10056
rect 7469 10047 7527 10053
rect 7469 10044 7481 10047
rect 7248 10016 7481 10044
rect 7248 10004 7254 10016
rect 7469 10013 7481 10016
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7561 10047 7619 10053
rect 7561 10013 7573 10047
rect 7607 10044 7619 10047
rect 7650 10044 7656 10056
rect 7607 10016 7656 10044
rect 7607 10013 7619 10016
rect 7561 10007 7619 10013
rect 7650 10004 7656 10016
rect 7708 10004 7714 10056
rect 10318 10004 10324 10056
rect 10376 10004 10382 10056
rect 10870 10004 10876 10056
rect 10928 10044 10934 10056
rect 12143 10047 12201 10053
rect 12143 10044 12155 10047
rect 10928 10016 12155 10044
rect 10928 10004 10934 10016
rect 12084 10013 12155 10016
rect 12189 10044 12201 10047
rect 12268 10044 12296 10084
rect 13740 10056 13768 10084
rect 14277 10081 14289 10115
rect 14323 10112 14335 10115
rect 15194 10112 15200 10124
rect 14323 10084 15200 10112
rect 14323 10081 14335 10084
rect 14277 10075 14335 10081
rect 15194 10072 15200 10084
rect 15252 10072 15258 10124
rect 16850 10072 16856 10124
rect 16908 10072 16914 10124
rect 13170 10044 13176 10056
rect 12189 10016 12296 10044
rect 12360 10016 13176 10044
rect 12189 10013 12204 10016
rect 12084 10012 12204 10013
rect 12143 10007 12201 10012
rect 6362 9976 6368 9988
rect 1688 9948 6368 9976
rect 6362 9936 6368 9948
rect 6420 9936 6426 9988
rect 11606 9936 11612 9988
rect 11664 9936 11670 9988
rect 11698 9936 11704 9988
rect 11756 9976 11762 9988
rect 11977 9979 12035 9985
rect 11977 9976 11989 9979
rect 11756 9948 11989 9976
rect 11756 9936 11762 9948
rect 11977 9945 11989 9948
rect 12023 9976 12035 9979
rect 12360 9976 12388 10016
rect 13170 10004 13176 10016
rect 13228 10004 13234 10056
rect 13265 10047 13323 10053
rect 13265 10013 13277 10047
rect 13311 10044 13323 10047
rect 13354 10044 13360 10056
rect 13311 10016 13360 10044
rect 13311 10013 13323 10016
rect 13265 10007 13323 10013
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 13446 10004 13452 10056
rect 13504 10044 13510 10056
rect 13504 10016 13676 10044
rect 13504 10004 13510 10016
rect 12023 9948 12388 9976
rect 12713 9979 12771 9985
rect 12023 9945 12035 9948
rect 11977 9939 12035 9945
rect 12713 9945 12725 9979
rect 12759 9976 12771 9979
rect 13648 9976 13676 10016
rect 13722 10004 13728 10056
rect 13780 10004 13786 10056
rect 13998 10044 14004 10056
rect 13832 10016 14004 10044
rect 13832 9976 13860 10016
rect 13998 10004 14004 10016
rect 14056 10044 14062 10056
rect 15473 10047 15531 10053
rect 15473 10044 15485 10047
rect 14056 10016 15485 10044
rect 14056 10004 14062 10016
rect 15473 10013 15485 10016
rect 15519 10013 15531 10047
rect 15473 10007 15531 10013
rect 15841 10047 15899 10053
rect 15841 10013 15853 10047
rect 15887 10044 15899 10047
rect 16666 10044 16672 10056
rect 15887 10016 16672 10044
rect 15887 10013 15899 10016
rect 15841 10007 15899 10013
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 12759 9948 13400 9976
rect 13648 9948 13860 9976
rect 14369 9979 14427 9985
rect 12759 9945 12771 9948
rect 12713 9939 12771 9945
rect 1854 9868 1860 9920
rect 1912 9868 1918 9920
rect 2682 9868 2688 9920
rect 2740 9868 2746 9920
rect 7742 9868 7748 9920
rect 7800 9868 7806 9920
rect 10413 9911 10471 9917
rect 10413 9877 10425 9911
rect 10459 9908 10471 9911
rect 10781 9911 10839 9917
rect 10781 9908 10793 9911
rect 10459 9880 10793 9908
rect 10459 9877 10471 9880
rect 10413 9871 10471 9877
rect 10781 9877 10793 9880
rect 10827 9877 10839 9911
rect 13372 9908 13400 9948
rect 14369 9945 14381 9979
rect 14415 9976 14427 9979
rect 14921 9979 14979 9985
rect 14921 9976 14933 9979
rect 14415 9948 14933 9976
rect 14415 9945 14427 9948
rect 14369 9939 14427 9945
rect 14921 9945 14933 9948
rect 14967 9945 14979 9979
rect 14921 9939 14979 9945
rect 13814 9908 13820 9920
rect 13372 9880 13820 9908
rect 10781 9871 10839 9877
rect 13814 9868 13820 9880
rect 13872 9868 13878 9920
rect 14458 9868 14464 9920
rect 14516 9868 14522 9920
rect 1104 9818 18124 9840
rect 1104 9766 3737 9818
rect 3789 9766 3801 9818
rect 3853 9766 3865 9818
rect 3917 9766 3929 9818
rect 3981 9766 3993 9818
rect 4045 9766 7992 9818
rect 8044 9766 8056 9818
rect 8108 9766 8120 9818
rect 8172 9766 8184 9818
rect 8236 9766 8248 9818
rect 8300 9766 12247 9818
rect 12299 9766 12311 9818
rect 12363 9766 12375 9818
rect 12427 9766 12439 9818
rect 12491 9766 12503 9818
rect 12555 9766 16502 9818
rect 16554 9766 16566 9818
rect 16618 9766 16630 9818
rect 16682 9766 16694 9818
rect 16746 9766 16758 9818
rect 16810 9766 18124 9818
rect 1104 9744 18124 9766
rect 2038 9664 2044 9716
rect 2096 9704 2102 9716
rect 7926 9704 7932 9716
rect 2096 9676 7932 9704
rect 2096 9664 2102 9676
rect 7926 9664 7932 9676
rect 7984 9664 7990 9716
rect 8864 9676 10548 9704
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 3016 9608 6224 9636
rect 3016 9596 3022 9608
rect 2225 9571 2283 9577
rect 2225 9537 2237 9571
rect 2271 9568 2283 9571
rect 2685 9571 2743 9577
rect 2685 9568 2697 9571
rect 2271 9540 2697 9568
rect 2271 9537 2283 9540
rect 2225 9531 2283 9537
rect 2685 9537 2697 9540
rect 2731 9537 2743 9571
rect 2685 9531 2743 9537
rect 3602 9528 3608 9580
rect 3660 9568 3666 9580
rect 3769 9571 3827 9577
rect 3769 9568 3781 9571
rect 3660 9540 3781 9568
rect 3660 9528 3666 9540
rect 3769 9537 3781 9540
rect 3815 9537 3827 9571
rect 3769 9531 3827 9537
rect 1673 9503 1731 9509
rect 1673 9469 1685 9503
rect 1719 9500 1731 9503
rect 2590 9500 2596 9512
rect 1719 9472 2596 9500
rect 1719 9469 1731 9472
rect 1673 9463 1731 9469
rect 2590 9460 2596 9472
rect 2648 9460 2654 9512
rect 2774 9460 2780 9512
rect 2832 9460 2838 9512
rect 2866 9460 2872 9512
rect 2924 9460 2930 9512
rect 3513 9503 3571 9509
rect 3513 9469 3525 9503
rect 3559 9469 3571 9503
rect 5537 9503 5595 9509
rect 5537 9500 5549 9503
rect 3513 9463 3571 9469
rect 4908 9472 5549 9500
rect 2130 9392 2136 9444
rect 2188 9432 2194 9444
rect 2188 9404 2774 9432
rect 2188 9392 2194 9404
rect 1762 9324 1768 9376
rect 1820 9364 1826 9376
rect 2317 9367 2375 9373
rect 2317 9364 2329 9367
rect 1820 9336 2329 9364
rect 1820 9324 1826 9336
rect 2317 9333 2329 9336
rect 2363 9333 2375 9367
rect 2746 9364 2774 9404
rect 3528 9364 3556 9463
rect 4706 9392 4712 9444
rect 4764 9432 4770 9444
rect 4908 9441 4936 9472
rect 5537 9469 5549 9472
rect 5583 9469 5595 9503
rect 6196 9500 6224 9608
rect 6362 9596 6368 9648
rect 6420 9596 6426 9648
rect 7558 9636 7564 9648
rect 6748 9608 7564 9636
rect 6270 9528 6276 9580
rect 6328 9568 6334 9580
rect 6549 9571 6607 9577
rect 6549 9568 6561 9571
rect 6328 9540 6561 9568
rect 6328 9528 6334 9540
rect 6549 9537 6561 9540
rect 6595 9537 6607 9571
rect 6549 9531 6607 9537
rect 6748 9500 6776 9608
rect 7558 9596 7564 9608
rect 7616 9636 7622 9648
rect 8864 9636 8892 9676
rect 7616 9608 8892 9636
rect 8956 9608 9444 9636
rect 7616 9596 7622 9608
rect 6932 9540 7788 9568
rect 6932 9512 6960 9540
rect 6196 9472 6776 9500
rect 6825 9503 6883 9509
rect 5537 9463 5595 9469
rect 6825 9469 6837 9503
rect 6871 9500 6883 9503
rect 6914 9500 6920 9512
rect 6871 9472 6920 9500
rect 6871 9469 6883 9472
rect 6825 9463 6883 9469
rect 6914 9460 6920 9472
rect 6972 9460 6978 9512
rect 7006 9460 7012 9512
rect 7064 9460 7070 9512
rect 7760 9500 7788 9540
rect 7834 9528 7840 9580
rect 7892 9568 7898 9580
rect 7929 9571 7987 9577
rect 7929 9568 7941 9571
rect 7892 9540 7941 9568
rect 7892 9528 7898 9540
rect 7929 9537 7941 9540
rect 7975 9537 7987 9571
rect 8570 9568 8576 9580
rect 7929 9531 7987 9537
rect 8128 9540 8576 9568
rect 8128 9500 8156 9540
rect 8570 9528 8576 9540
rect 8628 9528 8634 9580
rect 7760 9472 8156 9500
rect 8202 9460 8208 9512
rect 8260 9460 8266 9512
rect 8478 9460 8484 9512
rect 8536 9460 8542 9512
rect 8680 9500 8708 9608
rect 8846 9528 8852 9580
rect 8904 9568 8910 9580
rect 8956 9577 8984 9608
rect 8941 9571 8999 9577
rect 8941 9568 8953 9571
rect 8904 9540 8953 9568
rect 8904 9528 8910 9540
rect 8941 9537 8953 9540
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9568 9091 9571
rect 9122 9568 9128 9580
rect 9079 9540 9128 9568
rect 9079 9537 9091 9540
rect 9033 9531 9091 9537
rect 9122 9528 9128 9540
rect 9180 9528 9186 9580
rect 9416 9568 9444 9608
rect 9490 9596 9496 9648
rect 9548 9636 9554 9648
rect 10346 9639 10404 9645
rect 10346 9636 10358 9639
rect 9548 9608 10358 9636
rect 9548 9596 9554 9608
rect 10346 9605 10358 9608
rect 10392 9605 10404 9639
rect 10520 9636 10548 9676
rect 13262 9664 13268 9716
rect 13320 9664 13326 9716
rect 13446 9664 13452 9716
rect 13504 9664 13510 9716
rect 10520 9608 12434 9636
rect 10346 9599 10404 9605
rect 10229 9571 10287 9577
rect 10229 9568 10241 9571
rect 9416 9540 10241 9568
rect 10229 9537 10241 9540
rect 10275 9537 10287 9571
rect 10229 9531 10287 9537
rect 10778 9528 10784 9580
rect 10836 9528 10842 9580
rect 11422 9528 11428 9580
rect 11480 9568 11486 9580
rect 11609 9571 11667 9577
rect 11609 9568 11621 9571
rect 11480 9540 11621 9568
rect 11480 9528 11486 9540
rect 11609 9537 11621 9540
rect 11655 9537 11667 9571
rect 11609 9531 11667 9537
rect 11974 9528 11980 9580
rect 12032 9568 12038 9580
rect 12253 9571 12311 9577
rect 12253 9568 12265 9571
rect 12032 9540 12265 9568
rect 12032 9528 12038 9540
rect 12253 9537 12265 9540
rect 12299 9537 12311 9571
rect 12406 9568 12434 9608
rect 12802 9596 12808 9648
rect 12860 9636 12866 9648
rect 12989 9639 13047 9645
rect 12989 9636 13001 9639
rect 12860 9608 13001 9636
rect 12860 9596 12866 9608
rect 12989 9605 13001 9608
rect 13035 9605 13047 9639
rect 12989 9599 13047 9605
rect 14550 9596 14556 9648
rect 14608 9645 14614 9648
rect 14608 9636 14620 9645
rect 14608 9608 14653 9636
rect 14608 9599 14620 9608
rect 14608 9596 14614 9599
rect 15378 9568 15384 9580
rect 12406 9540 15384 9568
rect 12253 9531 12311 9537
rect 15378 9528 15384 9540
rect 15436 9528 15442 9580
rect 9401 9503 9459 9509
rect 9401 9500 9413 9503
rect 8680 9472 9413 9500
rect 9401 9469 9413 9472
rect 9447 9469 9459 9503
rect 9401 9463 9459 9469
rect 9493 9503 9551 9509
rect 9493 9469 9505 9503
rect 9539 9469 9551 9503
rect 9493 9463 9551 9469
rect 9861 9503 9919 9509
rect 9861 9469 9873 9503
rect 9907 9500 9919 9503
rect 10042 9500 10048 9512
rect 9907 9472 10048 9500
rect 9907 9469 9919 9472
rect 9861 9463 9919 9469
rect 4893 9435 4951 9441
rect 4893 9432 4905 9435
rect 4764 9404 4905 9432
rect 4764 9392 4770 9404
rect 4893 9401 4905 9404
rect 4939 9401 4951 9435
rect 4893 9395 4951 9401
rect 6178 9392 6184 9444
rect 6236 9432 6242 9444
rect 8113 9435 8171 9441
rect 8113 9432 8125 9435
rect 6236 9404 8125 9432
rect 6236 9392 6242 9404
rect 8113 9401 8125 9404
rect 8159 9401 8171 9435
rect 8220 9432 8248 9460
rect 9030 9432 9036 9444
rect 8220 9404 9036 9432
rect 8113 9395 8171 9401
rect 9030 9392 9036 9404
rect 9088 9392 9094 9444
rect 4154 9364 4160 9376
rect 2746 9336 4160 9364
rect 2317 9327 2375 9333
rect 4154 9324 4160 9336
rect 4212 9324 4218 9376
rect 4982 9324 4988 9376
rect 5040 9324 5046 9376
rect 6546 9324 6552 9376
rect 6604 9364 6610 9376
rect 6733 9367 6791 9373
rect 6733 9364 6745 9367
rect 6604 9336 6745 9364
rect 6604 9324 6610 9336
rect 6733 9333 6745 9336
rect 6779 9333 6791 9367
rect 6733 9327 6791 9333
rect 7190 9324 7196 9376
rect 7248 9364 7254 9376
rect 7653 9367 7711 9373
rect 7653 9364 7665 9367
rect 7248 9336 7665 9364
rect 7248 9324 7254 9336
rect 7653 9333 7665 9336
rect 7699 9333 7711 9367
rect 7653 9327 7711 9333
rect 7745 9367 7803 9373
rect 7745 9333 7757 9367
rect 7791 9364 7803 9367
rect 7926 9364 7932 9376
rect 7791 9336 7932 9364
rect 7791 9333 7803 9336
rect 7745 9327 7803 9333
rect 7926 9324 7932 9336
rect 7984 9324 7990 9376
rect 9508 9364 9536 9463
rect 10042 9460 10048 9472
rect 10100 9460 10106 9512
rect 10137 9503 10195 9509
rect 10137 9469 10149 9503
rect 10183 9469 10195 9503
rect 10137 9463 10195 9469
rect 10152 9432 10180 9463
rect 11238 9460 11244 9512
rect 11296 9500 11302 9512
rect 11882 9500 11888 9512
rect 11296 9472 11888 9500
rect 11296 9460 11302 9472
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 14829 9503 14887 9509
rect 14829 9469 14841 9503
rect 14875 9500 14887 9503
rect 15010 9500 15016 9512
rect 14875 9472 15016 9500
rect 14875 9469 14887 9472
rect 14829 9463 14887 9469
rect 15010 9460 15016 9472
rect 15068 9460 15074 9512
rect 15933 9503 15991 9509
rect 15933 9469 15945 9503
rect 15979 9500 15991 9503
rect 16298 9500 16304 9512
rect 15979 9472 16304 9500
rect 15979 9469 15991 9472
rect 15933 9463 15991 9469
rect 16298 9460 16304 9472
rect 16356 9460 16362 9512
rect 16390 9460 16396 9512
rect 16448 9500 16454 9512
rect 17221 9503 17279 9509
rect 17221 9500 17233 9503
rect 16448 9472 17233 9500
rect 16448 9460 16454 9472
rect 17221 9469 17233 9472
rect 17267 9469 17279 9503
rect 17221 9463 17279 9469
rect 10226 9432 10232 9444
rect 10152 9404 10232 9432
rect 10152 9364 10180 9404
rect 10226 9392 10232 9404
rect 10284 9392 10290 9444
rect 10505 9435 10563 9441
rect 10505 9401 10517 9435
rect 10551 9432 10563 9435
rect 11606 9432 11612 9444
rect 10551 9404 11612 9432
rect 10551 9401 10563 9404
rect 10505 9395 10563 9401
rect 11606 9392 11612 9404
rect 11664 9392 11670 9444
rect 15654 9392 15660 9444
rect 15712 9432 15718 9444
rect 16669 9435 16727 9441
rect 16669 9432 16681 9435
rect 15712 9404 16681 9432
rect 15712 9392 15718 9404
rect 16669 9401 16681 9404
rect 16715 9401 16727 9435
rect 16669 9395 16727 9401
rect 9508 9336 10180 9364
rect 10410 9324 10416 9376
rect 10468 9364 10474 9376
rect 10873 9367 10931 9373
rect 10873 9364 10885 9367
rect 10468 9336 10885 9364
rect 10468 9324 10474 9336
rect 10873 9333 10885 9336
rect 10919 9364 10931 9367
rect 11054 9364 11060 9376
rect 10919 9336 11060 9364
rect 10919 9333 10931 9336
rect 10873 9327 10931 9333
rect 11054 9324 11060 9336
rect 11112 9324 11118 9376
rect 12066 9324 12072 9376
rect 12124 9324 12130 9376
rect 16482 9324 16488 9376
rect 16540 9324 16546 9376
rect 1104 9274 18124 9296
rect 1104 9222 3077 9274
rect 3129 9222 3141 9274
rect 3193 9222 3205 9274
rect 3257 9222 3269 9274
rect 3321 9222 3333 9274
rect 3385 9222 7332 9274
rect 7384 9222 7396 9274
rect 7448 9222 7460 9274
rect 7512 9222 7524 9274
rect 7576 9222 7588 9274
rect 7640 9222 11587 9274
rect 11639 9222 11651 9274
rect 11703 9222 11715 9274
rect 11767 9222 11779 9274
rect 11831 9222 11843 9274
rect 11895 9222 15842 9274
rect 15894 9222 15906 9274
rect 15958 9222 15970 9274
rect 16022 9222 16034 9274
rect 16086 9222 16098 9274
rect 16150 9222 18124 9274
rect 1104 9200 18124 9222
rect 2866 9120 2872 9172
rect 2924 9160 2930 9172
rect 5166 9160 5172 9172
rect 2924 9132 5172 9160
rect 2924 9120 2930 9132
rect 5166 9120 5172 9132
rect 5224 9120 5230 9172
rect 6546 9120 6552 9172
rect 6604 9120 6610 9172
rect 6641 9163 6699 9169
rect 6641 9129 6653 9163
rect 6687 9160 6699 9163
rect 7006 9160 7012 9172
rect 6687 9132 7012 9160
rect 6687 9129 6699 9132
rect 6641 9123 6699 9129
rect 3513 9095 3571 9101
rect 3513 9061 3525 9095
rect 3559 9092 3571 9095
rect 4338 9092 4344 9104
rect 3559 9064 4344 9092
rect 3559 9061 3571 9064
rect 3513 9055 3571 9061
rect 4338 9052 4344 9064
rect 4396 9092 4402 9104
rect 4396 9064 5488 9092
rect 4396 9052 4402 9064
rect 4522 8984 4528 9036
rect 4580 8984 4586 9036
rect 4982 9024 4988 9036
rect 4632 8996 4988 9024
rect 1762 8916 1768 8968
rect 1820 8916 1826 8968
rect 1854 8916 1860 8968
rect 1912 8916 1918 8968
rect 2130 8916 2136 8968
rect 2188 8916 2194 8968
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8956 4307 8959
rect 4632 8956 4660 8996
rect 4982 8984 4988 8996
rect 5040 8984 5046 9036
rect 5258 8984 5264 9036
rect 5316 9024 5322 9036
rect 5353 9027 5411 9033
rect 5353 9024 5365 9027
rect 5316 8996 5365 9024
rect 5316 8984 5322 8996
rect 5353 8993 5365 8996
rect 5399 8993 5411 9027
rect 5460 9024 5488 9064
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 5460 8996 5641 9024
rect 5353 8987 5411 8993
rect 5629 8993 5641 8996
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 5902 8984 5908 9036
rect 5960 9024 5966 9036
rect 6086 9024 6092 9036
rect 5960 8996 6092 9024
rect 5960 8984 5966 8996
rect 6086 8984 6092 8996
rect 6144 8984 6150 9036
rect 4295 8928 4660 8956
rect 4295 8925 4307 8928
rect 4249 8919 4307 8925
rect 4706 8916 4712 8968
rect 4764 8916 4770 8968
rect 5810 8965 5816 8968
rect 4893 8959 4951 8965
rect 4893 8925 4905 8959
rect 4939 8925 4951 8959
rect 4893 8919 4951 8925
rect 5767 8959 5816 8965
rect 5767 8925 5779 8959
rect 5813 8925 5816 8959
rect 5767 8919 5816 8925
rect 2378 8891 2436 8897
rect 2378 8888 2390 8891
rect 2056 8860 2390 8888
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 1670 8820 1676 8832
rect 1627 8792 1676 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 1670 8780 1676 8792
rect 1728 8780 1734 8832
rect 2056 8829 2084 8860
rect 2378 8857 2390 8860
rect 2424 8857 2436 8891
rect 2378 8851 2436 8857
rect 2682 8848 2688 8900
rect 2740 8888 2746 8900
rect 3510 8888 3516 8900
rect 2740 8860 3516 8888
rect 2740 8848 2746 8860
rect 3510 8848 3516 8860
rect 3568 8888 3574 8900
rect 4341 8891 4399 8897
rect 4341 8888 4353 8891
rect 3568 8860 4353 8888
rect 3568 8848 3574 8860
rect 4341 8857 4353 8860
rect 4387 8888 4399 8891
rect 4614 8888 4620 8900
rect 4387 8860 4620 8888
rect 4387 8857 4399 8860
rect 4341 8851 4399 8857
rect 4614 8848 4620 8860
rect 4672 8848 4678 8900
rect 2041 8823 2099 8829
rect 2041 8789 2053 8823
rect 2087 8789 2099 8823
rect 2041 8783 2099 8789
rect 3881 8823 3939 8829
rect 3881 8789 3893 8823
rect 3927 8820 3939 8823
rect 4062 8820 4068 8832
rect 3927 8792 4068 8820
rect 3927 8789 3939 8792
rect 3881 8783 3939 8789
rect 4062 8780 4068 8792
rect 4120 8780 4126 8832
rect 4522 8780 4528 8832
rect 4580 8820 4586 8832
rect 4908 8820 4936 8919
rect 5810 8916 5816 8919
rect 5868 8916 5874 8968
rect 6656 8820 6684 9123
rect 7006 9120 7012 9132
rect 7064 9120 7070 9172
rect 7282 9120 7288 9172
rect 7340 9160 7346 9172
rect 8202 9160 8208 9172
rect 7340 9132 8208 9160
rect 7340 9120 7346 9132
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8665 9163 8723 9169
rect 8665 9129 8677 9163
rect 8711 9160 8723 9163
rect 9122 9160 9128 9172
rect 8711 9132 9128 9160
rect 8711 9129 8723 9132
rect 8665 9123 8723 9129
rect 9122 9120 9128 9132
rect 9180 9160 9186 9172
rect 10042 9160 10048 9172
rect 9180 9132 10048 9160
rect 9180 9120 9186 9132
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 10778 9120 10784 9172
rect 10836 9120 10842 9172
rect 11422 9120 11428 9172
rect 11480 9120 11486 9172
rect 12618 9120 12624 9172
rect 12676 9160 12682 9172
rect 13354 9160 13360 9172
rect 12676 9132 13360 9160
rect 12676 9120 12682 9132
rect 13354 9120 13360 9132
rect 13412 9120 13418 9172
rect 14277 9163 14335 9169
rect 14277 9129 14289 9163
rect 14323 9129 14335 9163
rect 14277 9123 14335 9129
rect 10226 9092 10232 9104
rect 9048 9064 10232 9092
rect 9048 9033 9076 9064
rect 10226 9052 10232 9064
rect 10284 9052 10290 9104
rect 13081 9095 13139 9101
rect 13081 9061 13093 9095
rect 13127 9061 13139 9095
rect 13081 9055 13139 9061
rect 8481 9027 8539 9033
rect 8481 8993 8493 9027
rect 8527 9024 8539 9027
rect 9033 9027 9091 9033
rect 9033 9024 9045 9027
rect 8527 8996 9045 9024
rect 8527 8993 8539 8996
rect 8481 8987 8539 8993
rect 9033 8993 9045 8996
rect 9079 8993 9091 9027
rect 10505 9027 10563 9033
rect 10505 9024 10517 9027
rect 9033 8987 9091 8993
rect 9508 8996 10517 9024
rect 9508 8968 9536 8996
rect 10505 8993 10517 8996
rect 10551 9024 10563 9027
rect 10873 9027 10931 9033
rect 10873 9024 10885 9027
rect 10551 8996 10885 9024
rect 10551 8993 10563 8996
rect 10505 8987 10563 8993
rect 10873 8993 10885 8996
rect 10919 8993 10931 9027
rect 10873 8987 10931 8993
rect 12986 8984 12992 9036
rect 13044 9024 13050 9036
rect 13096 9024 13124 9055
rect 13817 9027 13875 9033
rect 13817 9024 13829 9027
rect 13044 8996 13829 9024
rect 13044 8984 13050 8996
rect 13817 8993 13829 8996
rect 13863 9024 13875 9027
rect 14292 9024 14320 9123
rect 14550 9120 14556 9172
rect 14608 9160 14614 9172
rect 16390 9160 16396 9172
rect 14608 9132 16396 9160
rect 14608 9120 14614 9132
rect 16390 9120 16396 9132
rect 16448 9120 16454 9172
rect 14921 9095 14979 9101
rect 14921 9061 14933 9095
rect 14967 9061 14979 9095
rect 14921 9055 14979 9061
rect 13863 8996 14320 9024
rect 13863 8993 13875 8996
rect 13817 8987 13875 8993
rect 7742 8916 7748 8968
rect 7800 8965 7806 8968
rect 7800 8956 7812 8965
rect 7800 8928 7845 8956
rect 7800 8919 7812 8928
rect 7800 8916 7806 8919
rect 7926 8916 7932 8968
rect 7984 8956 7990 8968
rect 8021 8959 8079 8965
rect 8021 8956 8033 8959
rect 7984 8928 8033 8956
rect 7984 8916 7990 8928
rect 8021 8925 8033 8928
rect 8067 8925 8079 8959
rect 8021 8919 8079 8925
rect 8297 8959 8355 8965
rect 8297 8925 8309 8959
rect 8343 8925 8355 8959
rect 9490 8956 9496 8968
rect 8297 8919 8355 8925
rect 8496 8928 9496 8956
rect 8312 8888 8340 8919
rect 8496 8900 8524 8928
rect 9490 8916 9496 8928
rect 9548 8916 9554 8968
rect 10042 8916 10048 8968
rect 10100 8916 10106 8968
rect 10137 8959 10195 8965
rect 10137 8925 10149 8959
rect 10183 8956 10195 8959
rect 10226 8956 10232 8968
rect 10183 8928 10232 8956
rect 10183 8925 10195 8928
rect 10137 8919 10195 8925
rect 10226 8916 10232 8928
rect 10284 8916 10290 8968
rect 11241 8959 11299 8965
rect 11241 8956 11253 8959
rect 10428 8928 11253 8956
rect 8478 8888 8484 8900
rect 8312 8860 8484 8888
rect 8478 8848 8484 8860
rect 8536 8848 8542 8900
rect 8757 8891 8815 8897
rect 8757 8857 8769 8891
rect 8803 8888 8815 8891
rect 8846 8888 8852 8900
rect 8803 8860 8852 8888
rect 8803 8857 8815 8860
rect 8757 8851 8815 8857
rect 8846 8848 8852 8860
rect 8904 8848 8910 8900
rect 9125 8891 9183 8897
rect 9125 8857 9137 8891
rect 9171 8888 9183 8891
rect 9171 8860 9352 8888
rect 9171 8857 9183 8860
rect 9125 8851 9183 8857
rect 4580 8792 6684 8820
rect 4580 8780 4586 8792
rect 7650 8780 7656 8832
rect 7708 8820 7714 8832
rect 8113 8823 8171 8829
rect 8113 8820 8125 8823
rect 7708 8792 8125 8820
rect 7708 8780 7714 8792
rect 8113 8789 8125 8792
rect 8159 8789 8171 8823
rect 9324 8820 9352 8860
rect 9398 8848 9404 8900
rect 9456 8888 9462 8900
rect 10428 8897 10456 8928
rect 11241 8925 11253 8928
rect 11287 8925 11299 8959
rect 11241 8919 11299 8925
rect 11701 8959 11759 8965
rect 11701 8925 11713 8959
rect 11747 8956 11759 8959
rect 11747 8928 12434 8956
rect 11747 8925 11759 8928
rect 11701 8919 11759 8925
rect 9585 8891 9643 8897
rect 9585 8888 9597 8891
rect 9456 8860 9597 8888
rect 9456 8848 9462 8860
rect 9585 8857 9597 8860
rect 9631 8888 9643 8891
rect 10413 8891 10471 8897
rect 10413 8888 10425 8891
rect 9631 8860 10425 8888
rect 9631 8857 9643 8860
rect 9585 8851 9643 8857
rect 10413 8857 10425 8860
rect 10459 8857 10471 8891
rect 10413 8851 10471 8857
rect 10622 8891 10680 8897
rect 10622 8857 10634 8891
rect 10668 8888 10680 8891
rect 11968 8891 12026 8897
rect 10668 8860 10916 8888
rect 10668 8857 10680 8860
rect 10622 8851 10680 8857
rect 10888 8832 10916 8860
rect 11968 8857 11980 8891
rect 12014 8888 12026 8891
rect 12066 8888 12072 8900
rect 12014 8860 12072 8888
rect 12014 8857 12026 8860
rect 11968 8851 12026 8857
rect 12066 8848 12072 8860
rect 12124 8848 12130 8900
rect 12406 8888 12434 8928
rect 14366 8916 14372 8968
rect 14424 8956 14430 8968
rect 14553 8959 14611 8965
rect 14553 8956 14565 8959
rect 14424 8928 14565 8956
rect 14424 8916 14430 8928
rect 14553 8925 14565 8928
rect 14599 8925 14611 8959
rect 14553 8919 14611 8925
rect 12618 8888 12624 8900
rect 12406 8860 12624 8888
rect 12618 8848 12624 8860
rect 12676 8848 12682 8900
rect 13630 8848 13636 8900
rect 13688 8888 13694 8900
rect 14568 8888 14596 8919
rect 14734 8916 14740 8968
rect 14792 8916 14798 8968
rect 14826 8888 14832 8900
rect 13688 8860 14228 8888
rect 14568 8860 14832 8888
rect 13688 8848 13694 8860
rect 9674 8820 9680 8832
rect 9324 8792 9680 8820
rect 8113 8783 8171 8789
rect 9674 8780 9680 8792
rect 9732 8820 9738 8832
rect 10502 8820 10508 8832
rect 9732 8792 10508 8820
rect 9732 8780 9738 8792
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 10870 8780 10876 8832
rect 10928 8820 10934 8832
rect 11057 8823 11115 8829
rect 11057 8820 11069 8823
rect 10928 8792 11069 8820
rect 10928 8780 10934 8792
rect 11057 8789 11069 8792
rect 11103 8789 11115 8823
rect 11057 8783 11115 8789
rect 11146 8780 11152 8832
rect 11204 8820 11210 8832
rect 11882 8820 11888 8832
rect 11204 8792 11888 8820
rect 11204 8780 11210 8792
rect 11882 8780 11888 8792
rect 11940 8780 11946 8832
rect 13170 8780 13176 8832
rect 13228 8780 13234 8832
rect 13538 8780 13544 8832
rect 13596 8820 13602 8832
rect 14093 8823 14151 8829
rect 14093 8820 14105 8823
rect 13596 8792 14105 8820
rect 13596 8780 13602 8792
rect 14093 8789 14105 8792
rect 14139 8789 14151 8823
rect 14200 8820 14228 8860
rect 14826 8848 14832 8860
rect 14884 8848 14890 8900
rect 14936 8888 14964 9055
rect 16577 9027 16635 9033
rect 16577 9024 16589 9027
rect 16040 8996 16589 9024
rect 15010 8916 15016 8968
rect 15068 8916 15074 8968
rect 16040 8956 16068 8996
rect 16577 8993 16589 8996
rect 16623 9024 16635 9027
rect 17218 9024 17224 9036
rect 16623 8996 17224 9024
rect 16623 8993 16635 8996
rect 16577 8987 16635 8993
rect 17218 8984 17224 8996
rect 17276 8984 17282 9036
rect 15396 8928 16068 8956
rect 15396 8900 15424 8928
rect 16482 8916 16488 8968
rect 16540 8956 16546 8968
rect 16853 8959 16911 8965
rect 16853 8956 16865 8959
rect 16540 8928 16865 8956
rect 16540 8916 16546 8928
rect 16853 8925 16865 8928
rect 16899 8925 16911 8959
rect 17313 8959 17371 8965
rect 17313 8956 17325 8959
rect 16853 8919 16911 8925
rect 17236 8928 17325 8956
rect 15258 8891 15316 8897
rect 15258 8888 15270 8891
rect 14936 8860 15270 8888
rect 15258 8857 15270 8860
rect 15304 8857 15316 8891
rect 15258 8851 15316 8857
rect 15378 8848 15384 8900
rect 15436 8848 15442 8900
rect 15746 8888 15752 8900
rect 15488 8860 15752 8888
rect 15488 8820 15516 8860
rect 15746 8848 15752 8860
rect 15804 8848 15810 8900
rect 14200 8792 15516 8820
rect 14093 8783 14151 8789
rect 15562 8780 15568 8832
rect 15620 8820 15626 8832
rect 17236 8829 17264 8928
rect 17313 8925 17325 8928
rect 17359 8925 17371 8959
rect 17313 8919 17371 8925
rect 16761 8823 16819 8829
rect 16761 8820 16773 8823
rect 15620 8792 16773 8820
rect 15620 8780 15626 8792
rect 16761 8789 16773 8792
rect 16807 8789 16819 8823
rect 16761 8783 16819 8789
rect 17221 8823 17279 8829
rect 17221 8789 17233 8823
rect 17267 8789 17279 8823
rect 17221 8783 17279 8789
rect 17494 8780 17500 8832
rect 17552 8780 17558 8832
rect 1104 8730 18124 8752
rect 1104 8678 3737 8730
rect 3789 8678 3801 8730
rect 3853 8678 3865 8730
rect 3917 8678 3929 8730
rect 3981 8678 3993 8730
rect 4045 8678 7992 8730
rect 8044 8678 8056 8730
rect 8108 8678 8120 8730
rect 8172 8678 8184 8730
rect 8236 8678 8248 8730
rect 8300 8678 12247 8730
rect 12299 8678 12311 8730
rect 12363 8678 12375 8730
rect 12427 8678 12439 8730
rect 12491 8678 12503 8730
rect 12555 8678 16502 8730
rect 16554 8678 16566 8730
rect 16618 8678 16630 8730
rect 16682 8678 16694 8730
rect 16746 8678 16758 8730
rect 16810 8678 18124 8730
rect 1104 8656 18124 8678
rect 1854 8576 1860 8628
rect 1912 8616 1918 8628
rect 2961 8619 3019 8625
rect 2961 8616 2973 8619
rect 1912 8588 2973 8616
rect 1912 8576 1918 8588
rect 2961 8585 2973 8588
rect 3007 8585 3019 8619
rect 2961 8579 3019 8585
rect 3421 8619 3479 8625
rect 3421 8585 3433 8619
rect 3467 8616 3479 8619
rect 3510 8616 3516 8628
rect 3467 8588 3516 8616
rect 3467 8585 3479 8588
rect 3421 8579 3479 8585
rect 3510 8576 3516 8588
rect 3568 8576 3574 8628
rect 3602 8576 3608 8628
rect 3660 8616 3666 8628
rect 3973 8619 4031 8625
rect 3973 8616 3985 8619
rect 3660 8588 3985 8616
rect 3660 8576 3666 8588
rect 3973 8585 3985 8588
rect 4019 8585 4031 8619
rect 5350 8616 5356 8628
rect 3973 8579 4031 8585
rect 4540 8588 5356 8616
rect 2130 8548 2136 8560
rect 1412 8520 2136 8548
rect 1412 8489 1440 8520
rect 2130 8508 2136 8520
rect 2188 8508 2194 8560
rect 2590 8508 2596 8560
rect 2648 8548 2654 8560
rect 4540 8548 4568 8588
rect 5350 8576 5356 8588
rect 5408 8616 5414 8628
rect 5810 8616 5816 8628
rect 5408 8588 5816 8616
rect 5408 8576 5414 8588
rect 5810 8576 5816 8588
rect 5868 8576 5874 8628
rect 6178 8576 6184 8628
rect 6236 8576 6242 8628
rect 7190 8576 7196 8628
rect 7248 8616 7254 8628
rect 7285 8619 7343 8625
rect 7285 8616 7297 8619
rect 7248 8588 7297 8616
rect 7248 8576 7254 8588
rect 7285 8585 7297 8588
rect 7331 8585 7343 8619
rect 7285 8579 7343 8585
rect 7742 8576 7748 8628
rect 7800 8616 7806 8628
rect 8386 8616 8392 8628
rect 7800 8588 8392 8616
rect 7800 8576 7806 8588
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 9674 8616 9680 8628
rect 8588 8588 9680 8616
rect 2648 8520 4568 8548
rect 2648 8508 2654 8520
rect 7650 8508 7656 8560
rect 7708 8548 7714 8560
rect 8113 8551 8171 8557
rect 8113 8548 8125 8551
rect 7708 8520 8125 8548
rect 7708 8508 7714 8520
rect 8113 8517 8125 8520
rect 8159 8517 8171 8551
rect 8113 8511 8171 8517
rect 1670 8489 1676 8492
rect 1397 8483 1455 8489
rect 1397 8449 1409 8483
rect 1443 8449 1455 8483
rect 1664 8480 1676 8489
rect 1631 8452 1676 8480
rect 1397 8443 1455 8449
rect 1664 8443 1676 8452
rect 1670 8440 1676 8443
rect 1728 8440 1734 8492
rect 3329 8483 3387 8489
rect 3329 8449 3341 8483
rect 3375 8480 3387 8483
rect 3786 8480 3792 8492
rect 3375 8452 3792 8480
rect 3375 8449 3387 8452
rect 3329 8443 3387 8449
rect 3786 8440 3792 8452
rect 3844 8440 3850 8492
rect 4062 8440 4068 8492
rect 4120 8480 4126 8492
rect 4157 8483 4215 8489
rect 4157 8480 4169 8483
rect 4120 8452 4169 8480
rect 4120 8440 4126 8452
rect 4157 8449 4169 8452
rect 4203 8449 4215 8483
rect 4157 8443 4215 8449
rect 4341 8483 4399 8489
rect 4341 8449 4353 8483
rect 4387 8480 4399 8483
rect 4706 8480 4712 8492
rect 4387 8452 4712 8480
rect 4387 8449 4399 8452
rect 4341 8443 4399 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 5350 8440 5356 8492
rect 5408 8489 5414 8492
rect 5408 8483 5436 8489
rect 5424 8449 5436 8483
rect 5408 8443 5436 8449
rect 5408 8440 5414 8443
rect 7098 8440 7104 8492
rect 7156 8480 7162 8492
rect 7193 8483 7251 8489
rect 7193 8480 7205 8483
rect 7156 8452 7205 8480
rect 7156 8440 7162 8452
rect 7193 8449 7205 8452
rect 7239 8449 7251 8483
rect 7193 8443 7251 8449
rect 3602 8372 3608 8424
rect 3660 8372 3666 8424
rect 4522 8372 4528 8424
rect 4580 8372 4586 8424
rect 5261 8415 5319 8421
rect 5261 8412 5273 8415
rect 4724 8384 5273 8412
rect 2590 8304 2596 8356
rect 2648 8344 2654 8356
rect 2777 8347 2835 8353
rect 2777 8344 2789 8347
rect 2648 8316 2789 8344
rect 2648 8304 2654 8316
rect 2777 8313 2789 8316
rect 2823 8313 2835 8347
rect 2777 8307 2835 8313
rect 4338 8304 4344 8356
rect 4396 8344 4402 8356
rect 4724 8344 4752 8384
rect 5261 8381 5273 8384
rect 5307 8381 5319 8415
rect 5261 8375 5319 8381
rect 5537 8415 5595 8421
rect 5537 8381 5549 8415
rect 5583 8412 5595 8415
rect 5718 8412 5724 8424
rect 5583 8384 5724 8412
rect 5583 8381 5595 8384
rect 5537 8375 5595 8381
rect 5718 8372 5724 8384
rect 5776 8412 5782 8424
rect 6822 8412 6828 8424
rect 5776 8384 6828 8412
rect 5776 8372 5782 8384
rect 6822 8372 6828 8384
rect 6880 8372 6886 8424
rect 7009 8415 7067 8421
rect 7009 8381 7021 8415
rect 7055 8412 7067 8415
rect 8588 8412 8616 8588
rect 9674 8576 9680 8588
rect 9732 8576 9738 8628
rect 10505 8619 10563 8625
rect 10505 8585 10517 8619
rect 10551 8585 10563 8619
rect 10505 8579 10563 8585
rect 8662 8508 8668 8560
rect 8720 8548 8726 8560
rect 8757 8551 8815 8557
rect 8757 8548 8769 8551
rect 8720 8520 8769 8548
rect 8720 8508 8726 8520
rect 8757 8517 8769 8520
rect 8803 8548 8815 8551
rect 9030 8548 9036 8560
rect 8803 8520 9036 8548
rect 8803 8517 8815 8520
rect 8757 8511 8815 8517
rect 9030 8508 9036 8520
rect 9088 8508 9094 8560
rect 9217 8551 9275 8557
rect 9217 8517 9229 8551
rect 9263 8548 9275 8551
rect 10226 8548 10232 8560
rect 9263 8520 10232 8548
rect 9263 8517 9275 8520
rect 9217 8511 9275 8517
rect 10226 8508 10232 8520
rect 10284 8508 10290 8560
rect 10520 8548 10548 8579
rect 11974 8576 11980 8628
rect 12032 8576 12038 8628
rect 12345 8619 12403 8625
rect 12345 8585 12357 8619
rect 12391 8616 12403 8619
rect 13170 8616 13176 8628
rect 12391 8588 13176 8616
rect 12391 8585 12403 8588
rect 12345 8579 12403 8585
rect 13170 8576 13176 8588
rect 13228 8576 13234 8628
rect 13541 8619 13599 8625
rect 13541 8616 13553 8619
rect 13280 8588 13553 8616
rect 10781 8551 10839 8557
rect 10781 8548 10793 8551
rect 10520 8520 10793 8548
rect 10781 8517 10793 8520
rect 10827 8517 10839 8551
rect 10781 8511 10839 8517
rect 12437 8551 12495 8557
rect 12437 8517 12449 8551
rect 12483 8548 12495 8551
rect 12483 8520 12848 8548
rect 12483 8517 12495 8520
rect 12437 8511 12495 8517
rect 8846 8440 8852 8492
rect 8904 8480 8910 8492
rect 9125 8483 9183 8489
rect 9125 8480 9137 8483
rect 8904 8452 9137 8480
rect 8904 8440 8910 8452
rect 9125 8449 9137 8452
rect 9171 8480 9183 8483
rect 9398 8480 9404 8492
rect 9171 8452 9404 8480
rect 9171 8449 9183 8452
rect 9125 8443 9183 8449
rect 9398 8440 9404 8452
rect 9456 8440 9462 8492
rect 9490 8440 9496 8492
rect 9548 8480 9554 8492
rect 9677 8483 9735 8489
rect 9677 8480 9689 8483
rect 9548 8452 9689 8480
rect 9548 8440 9554 8452
rect 9677 8449 9689 8452
rect 9723 8480 9735 8483
rect 9861 8483 9919 8489
rect 9861 8480 9873 8483
rect 9723 8452 9873 8480
rect 9723 8449 9735 8452
rect 9677 8443 9735 8449
rect 9861 8449 9873 8452
rect 9907 8449 9919 8483
rect 10346 8483 10404 8489
rect 10346 8480 10358 8483
rect 9861 8443 9919 8449
rect 9968 8452 10358 8480
rect 7055 8384 8616 8412
rect 8665 8415 8723 8421
rect 7055 8381 7067 8384
rect 7009 8375 7067 8381
rect 7116 8356 7144 8384
rect 8665 8381 8677 8415
rect 8711 8381 8723 8415
rect 9416 8412 9444 8440
rect 9968 8412 9996 8452
rect 10346 8449 10358 8452
rect 10392 8449 10404 8483
rect 10346 8443 10404 8449
rect 11256 8452 12756 8480
rect 9416 8384 9996 8412
rect 8665 8375 8723 8381
rect 4396 8316 4752 8344
rect 4985 8347 5043 8353
rect 4396 8304 4402 8316
rect 4985 8313 4997 8347
rect 5031 8344 5043 8347
rect 5074 8344 5080 8356
rect 5031 8316 5080 8344
rect 5031 8313 5043 8316
rect 4985 8307 5043 8313
rect 5074 8304 5080 8316
rect 5132 8304 5138 8356
rect 7098 8304 7104 8356
rect 7156 8304 7162 8356
rect 7558 8304 7564 8356
rect 7616 8344 7622 8356
rect 7653 8347 7711 8353
rect 7653 8344 7665 8347
rect 7616 8316 7665 8344
rect 7616 8304 7622 8316
rect 7653 8313 7665 8316
rect 7699 8313 7711 8347
rect 8680 8344 8708 8375
rect 10042 8372 10048 8424
rect 10100 8412 10106 8424
rect 10137 8415 10195 8421
rect 10137 8412 10149 8415
rect 10100 8384 10149 8412
rect 10100 8372 10106 8384
rect 10137 8381 10149 8384
rect 10183 8381 10195 8415
rect 10137 8375 10195 8381
rect 10152 8344 10180 8375
rect 10226 8372 10232 8424
rect 10284 8412 10290 8424
rect 11146 8412 11152 8424
rect 10284 8384 11152 8412
rect 10284 8372 10290 8384
rect 11146 8372 11152 8384
rect 11204 8372 11210 8424
rect 10778 8344 10784 8356
rect 8680 8316 10784 8344
rect 7653 8307 7711 8313
rect 10778 8304 10784 8316
rect 10836 8304 10842 8356
rect 11256 8344 11284 8452
rect 12158 8372 12164 8424
rect 12216 8412 12222 8424
rect 12529 8415 12587 8421
rect 12529 8412 12541 8415
rect 12216 8384 12541 8412
rect 12216 8372 12222 8384
rect 12529 8381 12541 8384
rect 12575 8381 12587 8415
rect 12529 8375 12587 8381
rect 10888 8316 11284 8344
rect 12728 8344 12756 8452
rect 12820 8412 12848 8520
rect 12894 8508 12900 8560
rect 12952 8548 12958 8560
rect 13280 8548 13308 8588
rect 13541 8585 13553 8588
rect 13587 8616 13599 8619
rect 14274 8616 14280 8628
rect 13587 8588 14280 8616
rect 13587 8585 13599 8588
rect 13541 8579 13599 8585
rect 14274 8576 14280 8588
rect 14332 8576 14338 8628
rect 14734 8576 14740 8628
rect 14792 8616 14798 8628
rect 15197 8619 15255 8625
rect 15197 8616 15209 8619
rect 14792 8588 15209 8616
rect 14792 8576 14798 8588
rect 15197 8585 15209 8588
rect 15243 8585 15255 8619
rect 15197 8579 15255 8585
rect 15654 8576 15660 8628
rect 15712 8576 15718 8628
rect 15746 8576 15752 8628
rect 15804 8616 15810 8628
rect 17310 8616 17316 8628
rect 15804 8588 17316 8616
rect 15804 8576 15810 8588
rect 17310 8576 17316 8588
rect 17368 8576 17374 8628
rect 12952 8520 13308 8548
rect 12952 8508 12958 8520
rect 13446 8508 13452 8560
rect 13504 8548 13510 8560
rect 13722 8548 13728 8560
rect 13504 8520 13728 8548
rect 13504 8508 13510 8520
rect 13722 8508 13728 8520
rect 13780 8548 13786 8560
rect 13780 8520 17264 8548
rect 13780 8508 13786 8520
rect 13170 8440 13176 8492
rect 13228 8480 13234 8492
rect 13265 8483 13323 8489
rect 13265 8480 13277 8483
rect 13228 8452 13277 8480
rect 13228 8440 13234 8452
rect 13265 8449 13277 8452
rect 13311 8480 13323 8483
rect 13354 8480 13360 8492
rect 13311 8452 13360 8480
rect 13311 8449 13323 8452
rect 13265 8443 13323 8449
rect 13354 8440 13360 8452
rect 13412 8440 13418 8492
rect 13814 8440 13820 8492
rect 13872 8480 13878 8492
rect 14093 8483 14151 8489
rect 14093 8480 14105 8483
rect 13872 8452 14105 8480
rect 13872 8440 13878 8452
rect 14093 8449 14105 8452
rect 14139 8449 14151 8483
rect 14093 8443 14151 8449
rect 14108 8412 14136 8443
rect 14366 8440 14372 8492
rect 14424 8440 14430 8492
rect 14550 8440 14556 8492
rect 14608 8440 14614 8492
rect 15562 8480 15568 8492
rect 15028 8452 15568 8480
rect 14734 8412 14740 8424
rect 12820 8384 14044 8412
rect 14108 8384 14740 8412
rect 13630 8344 13636 8356
rect 12728 8316 13636 8344
rect 5092 8276 5120 8304
rect 6454 8276 6460 8288
rect 5092 8248 6460 8276
rect 6454 8236 6460 8248
rect 6512 8236 6518 8288
rect 8754 8236 8760 8288
rect 8812 8276 8818 8288
rect 9490 8276 9496 8288
rect 8812 8248 9496 8276
rect 8812 8236 8818 8248
rect 9490 8236 9496 8248
rect 9548 8276 9554 8288
rect 10888 8285 10916 8316
rect 13630 8304 13636 8316
rect 13688 8304 13694 8356
rect 14016 8344 14044 8384
rect 14734 8372 14740 8384
rect 14792 8372 14798 8424
rect 14016 8316 14320 8344
rect 10873 8279 10931 8285
rect 10873 8276 10885 8279
rect 9548 8248 10885 8276
rect 9548 8236 9554 8248
rect 10873 8245 10885 8248
rect 10919 8245 10931 8279
rect 10873 8239 10931 8245
rect 12066 8236 12072 8288
rect 12124 8276 12130 8288
rect 13814 8276 13820 8288
rect 12124 8248 13820 8276
rect 12124 8236 12130 8248
rect 13814 8236 13820 8248
rect 13872 8236 13878 8288
rect 13906 8236 13912 8288
rect 13964 8236 13970 8288
rect 14292 8276 14320 8316
rect 14366 8304 14372 8356
rect 14424 8344 14430 8356
rect 14918 8344 14924 8356
rect 14424 8316 14924 8344
rect 14424 8304 14430 8316
rect 14918 8304 14924 8316
rect 14976 8304 14982 8356
rect 15028 8276 15056 8452
rect 15562 8440 15568 8452
rect 15620 8440 15626 8492
rect 16206 8440 16212 8492
rect 16264 8480 16270 8492
rect 17236 8489 17264 8520
rect 16853 8483 16911 8489
rect 16853 8480 16865 8483
rect 16264 8452 16865 8480
rect 16264 8440 16270 8452
rect 16853 8449 16865 8452
rect 16899 8449 16911 8483
rect 16853 8443 16911 8449
rect 17221 8483 17279 8489
rect 17221 8449 17233 8483
rect 17267 8449 17279 8483
rect 17221 8443 17279 8449
rect 15194 8372 15200 8424
rect 15252 8412 15258 8424
rect 15470 8412 15476 8424
rect 15252 8384 15476 8412
rect 15252 8372 15258 8384
rect 15470 8372 15476 8384
rect 15528 8412 15534 8424
rect 15749 8415 15807 8421
rect 15749 8412 15761 8415
rect 15528 8384 15761 8412
rect 15528 8372 15534 8384
rect 15749 8381 15761 8384
rect 15795 8381 15807 8415
rect 15749 8375 15807 8381
rect 16301 8415 16359 8421
rect 16301 8381 16313 8415
rect 16347 8412 16359 8415
rect 16942 8412 16948 8424
rect 16347 8384 16948 8412
rect 16347 8381 16359 8384
rect 16301 8375 16359 8381
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 16390 8304 16396 8356
rect 16448 8344 16454 8356
rect 16669 8347 16727 8353
rect 16669 8344 16681 8347
rect 16448 8316 16681 8344
rect 16448 8304 16454 8316
rect 16669 8313 16681 8316
rect 16715 8313 16727 8347
rect 16669 8307 16727 8313
rect 14292 8248 15056 8276
rect 1104 8186 18124 8208
rect 1104 8134 3077 8186
rect 3129 8134 3141 8186
rect 3193 8134 3205 8186
rect 3257 8134 3269 8186
rect 3321 8134 3333 8186
rect 3385 8134 7332 8186
rect 7384 8134 7396 8186
rect 7448 8134 7460 8186
rect 7512 8134 7524 8186
rect 7576 8134 7588 8186
rect 7640 8134 11587 8186
rect 11639 8134 11651 8186
rect 11703 8134 11715 8186
rect 11767 8134 11779 8186
rect 11831 8134 11843 8186
rect 11895 8134 15842 8186
rect 15894 8134 15906 8186
rect 15958 8134 15970 8186
rect 16022 8134 16034 8186
rect 16086 8134 16098 8186
rect 16150 8134 18124 8186
rect 1104 8112 18124 8134
rect 3786 8032 3792 8084
rect 3844 8032 3850 8084
rect 10594 8032 10600 8084
rect 10652 8072 10658 8084
rect 10781 8075 10839 8081
rect 10781 8072 10793 8075
rect 10652 8044 10793 8072
rect 10652 8032 10658 8044
rect 10781 8041 10793 8044
rect 10827 8041 10839 8075
rect 10781 8035 10839 8041
rect 12345 8075 12403 8081
rect 12345 8041 12357 8075
rect 12391 8072 12403 8075
rect 12710 8072 12716 8084
rect 12391 8044 12716 8072
rect 12391 8041 12403 8044
rect 12345 8035 12403 8041
rect 4982 7964 4988 8016
rect 5040 8004 5046 8016
rect 5040 7976 7696 8004
rect 5040 7964 5046 7976
rect 4338 7896 4344 7948
rect 4396 7896 4402 7948
rect 7466 7936 7472 7948
rect 6932 7908 7472 7936
rect 5442 7828 5448 7880
rect 5500 7828 5506 7880
rect 5902 7828 5908 7880
rect 5960 7868 5966 7880
rect 6638 7868 6644 7880
rect 5960 7840 6644 7868
rect 5960 7828 5966 7840
rect 6638 7828 6644 7840
rect 6696 7868 6702 7880
rect 6932 7877 6960 7908
rect 7466 7896 7472 7908
rect 7524 7896 7530 7948
rect 7558 7896 7564 7948
rect 7616 7896 7622 7948
rect 7668 7936 7696 7976
rect 7742 7964 7748 8016
rect 7800 8004 7806 8016
rect 8205 8007 8263 8013
rect 8205 8004 8217 8007
rect 7800 7976 8217 8004
rect 7800 7964 7806 7976
rect 8205 7973 8217 7976
rect 8251 7973 8263 8007
rect 8205 7967 8263 7973
rect 7668 7908 7880 7936
rect 6917 7871 6975 7877
rect 6917 7868 6929 7871
rect 6696 7840 6929 7868
rect 6696 7828 6702 7840
rect 6917 7837 6929 7840
rect 6963 7837 6975 7871
rect 6917 7831 6975 7837
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7868 7435 7871
rect 7650 7868 7656 7880
rect 7423 7840 7656 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 4154 7760 4160 7812
rect 4212 7800 4218 7812
rect 4801 7803 4859 7809
rect 4801 7800 4813 7803
rect 4212 7772 4813 7800
rect 4212 7760 4218 7772
rect 4801 7769 4813 7772
rect 4847 7769 4859 7803
rect 4801 7763 4859 7769
rect 5534 7760 5540 7812
rect 5592 7800 5598 7812
rect 7208 7800 7236 7831
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 7852 7877 7880 7908
rect 7837 7871 7895 7877
rect 7837 7837 7849 7871
rect 7883 7837 7895 7871
rect 7837 7831 7895 7837
rect 10689 7871 10747 7877
rect 10689 7837 10701 7871
rect 10735 7868 10747 7871
rect 12360 7868 12388 8035
rect 12710 8032 12716 8044
rect 12768 8072 12774 8084
rect 12768 8044 12848 8072
rect 12768 8032 12774 8044
rect 12718 7881 12776 7887
rect 10735 7840 12388 7868
rect 10735 7837 10747 7840
rect 10689 7831 10747 7837
rect 10704 7800 10732 7831
rect 12526 7828 12532 7880
rect 12584 7828 12590 7880
rect 12718 7847 12730 7881
rect 12764 7878 12776 7881
rect 12820 7878 12848 8044
rect 12986 8032 12992 8084
rect 13044 8032 13050 8084
rect 16298 8032 16304 8084
rect 16356 8072 16362 8084
rect 16393 8075 16451 8081
rect 16393 8072 16405 8075
rect 16356 8044 16405 8072
rect 16356 8032 16362 8044
rect 16393 8041 16405 8044
rect 16439 8041 16451 8075
rect 16393 8035 16451 8041
rect 14550 7936 14556 7948
rect 13740 7908 14556 7936
rect 12764 7850 12848 7878
rect 12764 7847 12776 7850
rect 12718 7841 12776 7847
rect 13446 7828 13452 7880
rect 13504 7828 13510 7880
rect 13740 7877 13768 7908
rect 14550 7896 14556 7908
rect 14608 7896 14614 7948
rect 13725 7871 13783 7877
rect 13725 7837 13737 7871
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7868 13967 7871
rect 13998 7868 14004 7880
rect 13955 7840 14004 7868
rect 13955 7837 13967 7840
rect 13909 7831 13967 7837
rect 13998 7828 14004 7840
rect 14056 7828 14062 7880
rect 14366 7828 14372 7880
rect 14424 7828 14430 7880
rect 17773 7871 17831 7877
rect 17773 7868 17785 7871
rect 15672 7840 17785 7868
rect 5592 7772 10732 7800
rect 10980 7772 12434 7800
rect 5592 7760 5598 7772
rect 5258 7692 5264 7744
rect 5316 7692 5322 7744
rect 6546 7692 6552 7744
rect 6604 7732 6610 7744
rect 6733 7735 6791 7741
rect 6733 7732 6745 7735
rect 6604 7704 6745 7732
rect 6604 7692 6610 7704
rect 6733 7701 6745 7704
rect 6779 7701 6791 7735
rect 6733 7695 6791 7701
rect 7282 7692 7288 7744
rect 7340 7732 7346 7744
rect 7745 7735 7803 7741
rect 7745 7732 7757 7735
rect 7340 7704 7757 7732
rect 7340 7692 7346 7704
rect 7745 7701 7757 7704
rect 7791 7701 7803 7735
rect 7745 7695 7803 7701
rect 10318 7692 10324 7744
rect 10376 7732 10382 7744
rect 10980 7732 11008 7772
rect 10376 7704 11008 7732
rect 10376 7692 10382 7704
rect 11054 7692 11060 7744
rect 11112 7732 11118 7744
rect 11149 7735 11207 7741
rect 11149 7732 11161 7735
rect 11112 7704 11161 7732
rect 11112 7692 11118 7704
rect 11149 7701 11161 7704
rect 11195 7701 11207 7735
rect 12406 7732 12434 7772
rect 12802 7760 12808 7812
rect 12860 7800 12866 7812
rect 13265 7803 13323 7809
rect 13265 7800 13277 7803
rect 12860 7772 13277 7800
rect 12860 7760 12866 7772
rect 13265 7769 13277 7772
rect 13311 7769 13323 7803
rect 13265 7763 13323 7769
rect 12710 7732 12716 7744
rect 12406 7704 12716 7732
rect 11149 7695 11207 7701
rect 12710 7692 12716 7704
rect 12768 7692 12774 7744
rect 12986 7692 12992 7744
rect 13044 7732 13050 7744
rect 13173 7735 13231 7741
rect 13173 7732 13185 7735
rect 13044 7704 13185 7732
rect 13044 7692 13050 7704
rect 13173 7701 13185 7704
rect 13219 7701 13231 7735
rect 13173 7695 13231 7701
rect 14642 7692 14648 7744
rect 14700 7732 14706 7744
rect 15010 7732 15016 7744
rect 14700 7704 15016 7732
rect 14700 7692 14706 7704
rect 15010 7692 15016 7704
rect 15068 7732 15074 7744
rect 15672 7741 15700 7840
rect 17773 7837 17785 7840
rect 17819 7837 17831 7871
rect 17773 7831 17831 7837
rect 17494 7760 17500 7812
rect 17552 7809 17558 7812
rect 17552 7800 17564 7809
rect 17552 7772 17597 7800
rect 17552 7763 17564 7772
rect 17552 7760 17558 7763
rect 15657 7735 15715 7741
rect 15657 7732 15669 7735
rect 15068 7704 15669 7732
rect 15068 7692 15074 7704
rect 15657 7701 15669 7704
rect 15703 7701 15715 7735
rect 15657 7695 15715 7701
rect 1104 7642 18124 7664
rect 1104 7590 3737 7642
rect 3789 7590 3801 7642
rect 3853 7590 3865 7642
rect 3917 7590 3929 7642
rect 3981 7590 3993 7642
rect 4045 7590 7992 7642
rect 8044 7590 8056 7642
rect 8108 7590 8120 7642
rect 8172 7590 8184 7642
rect 8236 7590 8248 7642
rect 8300 7590 12247 7642
rect 12299 7590 12311 7642
rect 12363 7590 12375 7642
rect 12427 7590 12439 7642
rect 12491 7590 12503 7642
rect 12555 7590 16502 7642
rect 16554 7590 16566 7642
rect 16618 7590 16630 7642
rect 16682 7590 16694 7642
rect 16746 7590 16758 7642
rect 16810 7590 18124 7642
rect 1104 7568 18124 7590
rect 7282 7488 7288 7540
rect 7340 7488 7346 7540
rect 7466 7488 7472 7540
rect 7524 7528 7530 7540
rect 10318 7528 10324 7540
rect 7524 7500 10324 7528
rect 7524 7488 7530 7500
rect 10318 7488 10324 7500
rect 10376 7488 10382 7540
rect 12710 7488 12716 7540
rect 12768 7528 12774 7540
rect 13538 7528 13544 7540
rect 12768 7500 13544 7528
rect 12768 7488 12774 7500
rect 13538 7488 13544 7500
rect 13596 7488 13602 7540
rect 13817 7531 13875 7537
rect 13817 7497 13829 7531
rect 13863 7497 13875 7531
rect 13817 7491 13875 7497
rect 14185 7531 14243 7537
rect 14185 7497 14197 7531
rect 14231 7528 14243 7531
rect 14458 7528 14464 7540
rect 14231 7500 14464 7528
rect 14231 7497 14243 7500
rect 14185 7491 14243 7497
rect 3329 7463 3387 7469
rect 3329 7429 3341 7463
rect 3375 7460 3387 7463
rect 4982 7460 4988 7472
rect 3375 7432 4988 7460
rect 3375 7429 3387 7432
rect 3329 7423 3387 7429
rect 4982 7420 4988 7432
rect 5040 7420 5046 7472
rect 6181 7463 6239 7469
rect 6181 7429 6193 7463
rect 6227 7460 6239 7463
rect 7374 7460 7380 7472
rect 6227 7432 7380 7460
rect 6227 7429 6239 7432
rect 6181 7423 6239 7429
rect 7374 7420 7380 7432
rect 7432 7420 7438 7472
rect 9582 7420 9588 7472
rect 9640 7460 9646 7472
rect 10689 7463 10747 7469
rect 10689 7460 10701 7463
rect 9640 7432 10701 7460
rect 9640 7420 9646 7432
rect 10689 7429 10701 7432
rect 10735 7429 10747 7463
rect 12066 7460 12072 7472
rect 10689 7423 10747 7429
rect 11716 7432 12072 7460
rect 3237 7395 3295 7401
rect 3237 7361 3249 7395
rect 3283 7392 3295 7395
rect 3697 7395 3755 7401
rect 3697 7392 3709 7395
rect 3283 7364 3709 7392
rect 3283 7361 3295 7364
rect 3237 7355 3295 7361
rect 3697 7361 3709 7364
rect 3743 7361 3755 7395
rect 3697 7355 3755 7361
rect 4154 7352 4160 7404
rect 4212 7392 4218 7404
rect 4433 7395 4491 7401
rect 4433 7392 4445 7395
rect 4212 7364 4445 7392
rect 4212 7352 4218 7364
rect 4433 7361 4445 7364
rect 4479 7361 4491 7395
rect 4433 7355 4491 7361
rect 9122 7352 9128 7404
rect 9180 7392 9186 7404
rect 9473 7395 9531 7401
rect 9473 7392 9485 7395
rect 9180 7364 9485 7392
rect 9180 7352 9186 7364
rect 9473 7361 9485 7364
rect 9519 7361 9531 7395
rect 9473 7355 9531 7361
rect 9766 7352 9772 7404
rect 9824 7392 9830 7404
rect 11716 7401 11744 7432
rect 12066 7420 12072 7432
rect 12124 7420 12130 7472
rect 12986 7420 12992 7472
rect 13044 7460 13050 7472
rect 13449 7463 13507 7469
rect 13449 7460 13461 7463
rect 13044 7432 13461 7460
rect 13044 7420 13050 7432
rect 13449 7429 13461 7432
rect 13495 7429 13507 7463
rect 13449 7423 13507 7429
rect 11701 7395 11759 7401
rect 9824 7364 11376 7392
rect 9824 7352 9830 7364
rect 2958 7284 2964 7336
rect 3016 7324 3022 7336
rect 3421 7327 3479 7333
rect 3421 7324 3433 7327
rect 3016 7296 3433 7324
rect 3016 7284 3022 7296
rect 3421 7293 3433 7296
rect 3467 7293 3479 7327
rect 3421 7287 3479 7293
rect 4246 7284 4252 7336
rect 4304 7284 4310 7336
rect 6733 7327 6791 7333
rect 6733 7293 6745 7327
rect 6779 7324 6791 7327
rect 7650 7324 7656 7336
rect 6779 7296 7656 7324
rect 6779 7293 6791 7296
rect 6733 7287 6791 7293
rect 7650 7284 7656 7296
rect 7708 7284 7714 7336
rect 9217 7327 9275 7333
rect 9217 7324 9229 7327
rect 8680 7296 9229 7324
rect 2866 7148 2872 7200
rect 2924 7148 2930 7200
rect 8202 7148 8208 7200
rect 8260 7188 8266 7200
rect 8680 7197 8708 7296
rect 9217 7293 9229 7296
rect 9263 7293 9275 7327
rect 11241 7327 11299 7333
rect 11241 7324 11253 7327
rect 9217 7287 9275 7293
rect 10612 7296 11253 7324
rect 10612 7200 10640 7296
rect 11241 7293 11253 7296
rect 11287 7293 11299 7327
rect 11348 7324 11376 7364
rect 11701 7361 11713 7395
rect 11747 7361 11759 7395
rect 11701 7355 11759 7361
rect 11974 7352 11980 7404
rect 12032 7352 12038 7404
rect 12158 7352 12164 7404
rect 12216 7352 12222 7404
rect 12342 7352 12348 7404
rect 12400 7352 12406 7404
rect 12526 7401 12532 7404
rect 12493 7395 12532 7401
rect 12493 7361 12505 7395
rect 12493 7355 12532 7361
rect 12508 7352 12532 7355
rect 12584 7352 12590 7404
rect 12621 7395 12679 7401
rect 12621 7361 12633 7395
rect 12667 7361 12679 7395
rect 12621 7355 12679 7361
rect 12508 7324 12536 7352
rect 11348 7296 12536 7324
rect 12636 7324 12664 7355
rect 12710 7352 12716 7404
rect 12768 7352 12774 7404
rect 12802 7352 12808 7404
rect 12860 7401 12866 7404
rect 12860 7392 12868 7401
rect 12860 7364 12905 7392
rect 12860 7355 12868 7364
rect 12860 7352 12866 7355
rect 13078 7352 13084 7404
rect 13136 7352 13142 7404
rect 13262 7401 13268 7404
rect 13229 7395 13268 7401
rect 13229 7361 13241 7395
rect 13229 7355 13268 7361
rect 13262 7352 13268 7355
rect 13320 7352 13326 7404
rect 13630 7401 13636 7404
rect 13357 7395 13415 7401
rect 13357 7361 13369 7395
rect 13403 7361 13415 7395
rect 13357 7355 13415 7361
rect 13587 7395 13636 7401
rect 13587 7361 13599 7395
rect 13633 7361 13636 7395
rect 13587 7355 13636 7361
rect 12986 7324 12992 7336
rect 12636 7296 12992 7324
rect 11241 7287 11299 7293
rect 12986 7284 12992 7296
rect 13044 7284 13050 7336
rect 13372 7324 13400 7355
rect 13630 7352 13636 7355
rect 13688 7352 13694 7404
rect 13832 7324 13860 7491
rect 14458 7488 14464 7500
rect 14516 7528 14522 7540
rect 16298 7528 16304 7540
rect 14516 7500 16304 7528
rect 14516 7488 14522 7500
rect 16298 7488 16304 7500
rect 16356 7488 16362 7540
rect 13906 7420 13912 7472
rect 13964 7460 13970 7472
rect 13964 7432 16528 7460
rect 13964 7420 13970 7432
rect 13998 7352 14004 7404
rect 14056 7392 14062 7404
rect 15102 7392 15108 7404
rect 14056 7364 15108 7392
rect 14056 7352 14062 7364
rect 15102 7352 15108 7364
rect 15160 7352 15166 7404
rect 16229 7395 16287 7401
rect 16229 7361 16241 7395
rect 16275 7392 16287 7395
rect 16390 7392 16396 7404
rect 16275 7364 16396 7392
rect 16275 7361 16287 7364
rect 16229 7355 16287 7361
rect 16390 7352 16396 7364
rect 16448 7352 16454 7404
rect 16500 7401 16528 7432
rect 16485 7395 16543 7401
rect 16485 7361 16497 7395
rect 16531 7361 16543 7395
rect 16485 7355 16543 7361
rect 17770 7352 17776 7404
rect 17828 7352 17834 7404
rect 13372 7296 13860 7324
rect 14274 7284 14280 7336
rect 14332 7284 14338 7336
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7324 14519 7327
rect 14550 7324 14556 7336
rect 14507 7296 14556 7324
rect 14507 7293 14519 7296
rect 14461 7287 14519 7293
rect 14550 7284 14556 7296
rect 14608 7284 14614 7336
rect 14642 7284 14648 7336
rect 14700 7284 14706 7336
rect 17497 7327 17555 7333
rect 17497 7293 17509 7327
rect 17543 7293 17555 7327
rect 17497 7287 17555 7293
rect 12158 7216 12164 7268
rect 12216 7256 12222 7268
rect 15010 7256 15016 7268
rect 12216 7228 15016 7256
rect 12216 7216 12222 7228
rect 15010 7216 15016 7228
rect 15068 7256 15074 7268
rect 15105 7259 15163 7265
rect 15105 7256 15117 7259
rect 15068 7228 15117 7256
rect 15068 7216 15074 7228
rect 15105 7225 15117 7228
rect 15151 7225 15163 7259
rect 15105 7219 15163 7225
rect 8665 7191 8723 7197
rect 8665 7188 8677 7191
rect 8260 7160 8677 7188
rect 8260 7148 8266 7160
rect 8665 7157 8677 7160
rect 8711 7157 8723 7191
rect 8665 7151 8723 7157
rect 10594 7148 10600 7200
rect 10652 7148 10658 7200
rect 11146 7148 11152 7200
rect 11204 7188 11210 7200
rect 11517 7191 11575 7197
rect 11517 7188 11529 7191
rect 11204 7160 11529 7188
rect 11204 7148 11210 7160
rect 11517 7157 11529 7160
rect 11563 7157 11575 7191
rect 11517 7151 11575 7157
rect 12526 7148 12532 7200
rect 12584 7188 12590 7200
rect 12894 7188 12900 7200
rect 12584 7160 12900 7188
rect 12584 7148 12590 7160
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 12989 7191 13047 7197
rect 12989 7157 13001 7191
rect 13035 7188 13047 7191
rect 13630 7188 13636 7200
rect 13035 7160 13636 7188
rect 13035 7157 13047 7160
rect 12989 7151 13047 7157
rect 13630 7148 13636 7160
rect 13688 7148 13694 7200
rect 13725 7191 13783 7197
rect 13725 7157 13737 7191
rect 13771 7188 13783 7191
rect 14182 7188 14188 7200
rect 13771 7160 14188 7188
rect 13771 7157 13783 7160
rect 13725 7151 13783 7157
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 14734 7148 14740 7200
rect 14792 7188 14798 7200
rect 17512 7188 17540 7287
rect 14792 7160 17540 7188
rect 14792 7148 14798 7160
rect 1104 7098 18124 7120
rect 1104 7046 3077 7098
rect 3129 7046 3141 7098
rect 3193 7046 3205 7098
rect 3257 7046 3269 7098
rect 3321 7046 3333 7098
rect 3385 7046 7332 7098
rect 7384 7046 7396 7098
rect 7448 7046 7460 7098
rect 7512 7046 7524 7098
rect 7576 7046 7588 7098
rect 7640 7046 11587 7098
rect 11639 7046 11651 7098
rect 11703 7046 11715 7098
rect 11767 7046 11779 7098
rect 11831 7046 11843 7098
rect 11895 7046 15842 7098
rect 15894 7046 15906 7098
rect 15958 7046 15970 7098
rect 16022 7046 16034 7098
rect 16086 7046 16098 7098
rect 16150 7046 18124 7098
rect 1104 7024 18124 7046
rect 5537 6987 5595 6993
rect 5537 6953 5549 6987
rect 5583 6984 5595 6987
rect 6178 6984 6184 6996
rect 5583 6956 6184 6984
rect 5583 6953 5595 6956
rect 5537 6947 5595 6953
rect 6178 6944 6184 6956
rect 6236 6944 6242 6996
rect 7377 6987 7435 6993
rect 7377 6953 7389 6987
rect 7423 6984 7435 6987
rect 7650 6984 7656 6996
rect 7423 6956 7656 6984
rect 7423 6953 7435 6956
rect 7377 6947 7435 6953
rect 7650 6944 7656 6956
rect 7708 6944 7714 6996
rect 10229 6987 10287 6993
rect 7760 6956 9674 6984
rect 5994 6876 6000 6928
rect 6052 6876 6058 6928
rect 7760 6916 7788 6956
rect 7024 6888 7788 6916
rect 9646 6916 9674 6956
rect 10229 6953 10241 6987
rect 10275 6984 10287 6987
rect 10594 6984 10600 6996
rect 10275 6956 10600 6984
rect 10275 6953 10287 6956
rect 10229 6947 10287 6953
rect 10594 6944 10600 6956
rect 10652 6944 10658 6996
rect 12342 6984 12348 6996
rect 10704 6956 12348 6984
rect 10502 6916 10508 6928
rect 9646 6888 10508 6916
rect 6012 6848 6040 6876
rect 7024 6848 7052 6888
rect 10502 6876 10508 6888
rect 10560 6916 10566 6928
rect 10704 6916 10732 6956
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 12986 6944 12992 6996
rect 13044 6984 13050 6996
rect 14093 6987 14151 6993
rect 14093 6984 14105 6987
rect 13044 6956 14105 6984
rect 13044 6944 13050 6956
rect 14093 6953 14105 6956
rect 14139 6953 14151 6987
rect 14093 6947 14151 6953
rect 14826 6944 14832 6996
rect 14884 6984 14890 6996
rect 15013 6987 15071 6993
rect 15013 6984 15025 6987
rect 14884 6956 15025 6984
rect 14884 6944 14890 6956
rect 15013 6953 15025 6956
rect 15059 6953 15071 6987
rect 15013 6947 15071 6953
rect 10560 6888 10732 6916
rect 10560 6876 10566 6888
rect 14734 6876 14740 6928
rect 14792 6916 14798 6928
rect 14792 6888 16436 6916
rect 14792 6876 14798 6888
rect 7650 6848 7656 6860
rect 5920 6820 7052 6848
rect 7116 6820 7656 6848
rect 2041 6783 2099 6789
rect 2041 6749 2053 6783
rect 2087 6780 2099 6783
rect 4154 6780 4160 6792
rect 2087 6752 4160 6780
rect 2087 6749 2099 6752
rect 2041 6743 2099 6749
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 4424 6783 4482 6789
rect 4424 6749 4436 6783
rect 4470 6780 4482 6783
rect 5258 6780 5264 6792
rect 4470 6752 5264 6780
rect 4470 6749 4482 6752
rect 4424 6743 4482 6749
rect 5258 6740 5264 6752
rect 5316 6740 5322 6792
rect 5920 6789 5948 6820
rect 6086 6789 6092 6792
rect 5905 6783 5963 6789
rect 5905 6749 5917 6783
rect 5951 6749 5963 6783
rect 5905 6743 5963 6749
rect 6053 6783 6092 6789
rect 6053 6749 6065 6783
rect 6053 6743 6092 6749
rect 6086 6740 6092 6743
rect 6144 6740 6150 6792
rect 7116 6789 7144 6820
rect 7650 6808 7656 6820
rect 7708 6808 7714 6860
rect 9030 6808 9036 6860
rect 9088 6848 9094 6860
rect 9677 6851 9735 6857
rect 9677 6848 9689 6851
rect 9088 6820 9689 6848
rect 9088 6808 9094 6820
rect 9677 6817 9689 6820
rect 9723 6817 9735 6851
rect 12158 6848 12164 6860
rect 9677 6811 9735 6817
rect 11716 6820 12164 6848
rect 6411 6783 6469 6789
rect 6411 6749 6423 6783
rect 6457 6780 6469 6783
rect 6641 6783 6699 6789
rect 6641 6780 6653 6783
rect 6457 6752 6653 6780
rect 6457 6749 6469 6752
rect 6411 6743 6469 6749
rect 6641 6749 6653 6752
rect 6687 6749 6699 6783
rect 6641 6743 6699 6749
rect 6825 6783 6883 6789
rect 6825 6749 6837 6783
rect 6871 6749 6883 6783
rect 6825 6743 6883 6749
rect 7101 6783 7159 6789
rect 7101 6749 7113 6783
rect 7147 6749 7159 6783
rect 7101 6743 7159 6749
rect 7285 6783 7343 6789
rect 7285 6749 7297 6783
rect 7331 6780 7343 6783
rect 8202 6780 8208 6792
rect 7331 6752 7788 6780
rect 7331 6749 7343 6752
rect 7285 6743 7343 6749
rect 2308 6715 2366 6721
rect 2308 6681 2320 6715
rect 2354 6712 2366 6715
rect 2498 6712 2504 6724
rect 2354 6684 2504 6712
rect 2354 6681 2366 6684
rect 2308 6675 2366 6681
rect 2498 6672 2504 6684
rect 2556 6672 2562 6724
rect 4522 6672 4528 6724
rect 4580 6712 4586 6724
rect 6181 6715 6239 6721
rect 6181 6712 6193 6715
rect 4580 6684 6193 6712
rect 4580 6672 4586 6684
rect 6181 6681 6193 6684
rect 6227 6681 6239 6715
rect 6181 6675 6239 6681
rect 6273 6715 6331 6721
rect 6273 6681 6285 6715
rect 6319 6712 6331 6715
rect 6730 6712 6736 6724
rect 6319 6684 6736 6712
rect 6319 6681 6331 6684
rect 6273 6675 6331 6681
rect 6730 6672 6736 6684
rect 6788 6672 6794 6724
rect 6840 6712 6868 6743
rect 7650 6712 7656 6724
rect 6840 6684 7656 6712
rect 7650 6672 7656 6684
rect 7708 6672 7714 6724
rect 3421 6647 3479 6653
rect 3421 6613 3433 6647
rect 3467 6644 3479 6647
rect 4246 6644 4252 6656
rect 3467 6616 4252 6644
rect 3467 6613 3479 6616
rect 3421 6607 3479 6613
rect 4246 6604 4252 6616
rect 4304 6604 4310 6656
rect 6549 6647 6607 6653
rect 6549 6613 6561 6647
rect 6595 6644 6607 6647
rect 6822 6644 6828 6656
rect 6595 6616 6828 6644
rect 6595 6613 6607 6616
rect 6549 6607 6607 6613
rect 6822 6604 6828 6616
rect 6880 6604 6886 6656
rect 7558 6604 7564 6656
rect 7616 6644 7622 6656
rect 7760 6644 7788 6752
rect 7852 6752 8208 6780
rect 7852 6724 7880 6752
rect 8202 6740 8208 6752
rect 8260 6780 8266 6792
rect 8757 6783 8815 6789
rect 8757 6780 8769 6783
rect 8260 6752 8769 6780
rect 8260 6740 8266 6752
rect 8757 6749 8769 6752
rect 8803 6749 8815 6783
rect 8757 6743 8815 6749
rect 9493 6783 9551 6789
rect 9493 6749 9505 6783
rect 9539 6780 9551 6783
rect 9582 6780 9588 6792
rect 9539 6752 9588 6780
rect 9539 6749 9551 6752
rect 9493 6743 9551 6749
rect 9582 6740 9588 6752
rect 9640 6740 9646 6792
rect 9950 6740 9956 6792
rect 10008 6740 10014 6792
rect 10502 6740 10508 6792
rect 10560 6740 10566 6792
rect 11716 6789 11744 6820
rect 12158 6808 12164 6820
rect 12216 6808 12222 6860
rect 14090 6808 14096 6860
rect 14148 6848 14154 6860
rect 14645 6851 14703 6857
rect 14645 6848 14657 6851
rect 14148 6820 14657 6848
rect 14148 6808 14154 6820
rect 14645 6817 14657 6820
rect 14691 6817 14703 6851
rect 14645 6811 14703 6817
rect 10598 6783 10656 6789
rect 10598 6749 10610 6783
rect 10644 6749 10656 6783
rect 10598 6743 10656 6749
rect 11009 6783 11067 6789
rect 11009 6749 11021 6783
rect 11055 6780 11067 6783
rect 11241 6783 11299 6789
rect 11241 6780 11253 6783
rect 11055 6752 11253 6780
rect 11055 6749 11067 6752
rect 11009 6743 11067 6749
rect 11241 6749 11253 6752
rect 11287 6749 11299 6783
rect 11241 6743 11299 6749
rect 11425 6783 11483 6789
rect 11425 6749 11437 6783
rect 11471 6749 11483 6783
rect 11425 6743 11483 6749
rect 11701 6783 11759 6789
rect 11701 6749 11713 6783
rect 11747 6749 11759 6783
rect 11701 6743 11759 6749
rect 7834 6672 7840 6724
rect 7892 6672 7898 6724
rect 8386 6672 8392 6724
rect 8444 6712 8450 6724
rect 8490 6715 8548 6721
rect 8490 6712 8502 6715
rect 8444 6684 8502 6712
rect 8444 6672 8450 6684
rect 8490 6681 8502 6684
rect 8536 6681 8548 6715
rect 9968 6712 9996 6740
rect 10612 6712 10640 6743
rect 8490 6675 8548 6681
rect 8588 6684 9996 6712
rect 10336 6684 10640 6712
rect 8588 6644 8616 6684
rect 7616 6616 8616 6644
rect 7616 6604 7622 6616
rect 8938 6604 8944 6656
rect 8996 6644 9002 6656
rect 9125 6647 9183 6653
rect 9125 6644 9137 6647
rect 8996 6616 9137 6644
rect 8996 6604 9002 6616
rect 9125 6613 9137 6616
rect 9171 6613 9183 6647
rect 9125 6607 9183 6613
rect 9582 6604 9588 6656
rect 9640 6604 9646 6656
rect 9766 6604 9772 6656
rect 9824 6644 9830 6656
rect 10336 6644 10364 6684
rect 10778 6672 10784 6724
rect 10836 6672 10842 6724
rect 10873 6715 10931 6721
rect 10873 6681 10885 6715
rect 10919 6681 10931 6715
rect 11440 6712 11468 6743
rect 11882 6740 11888 6792
rect 11940 6740 11946 6792
rect 13909 6783 13967 6789
rect 13909 6749 13921 6783
rect 13955 6780 13967 6783
rect 14366 6780 14372 6792
rect 13955 6752 14372 6780
rect 13955 6749 13967 6752
rect 13909 6743 13967 6749
rect 14366 6740 14372 6752
rect 14424 6740 14430 6792
rect 14458 6740 14464 6792
rect 14516 6740 14522 6792
rect 14660 6780 14688 6811
rect 15470 6808 15476 6860
rect 15528 6808 15534 6860
rect 16408 6857 16436 6888
rect 16393 6851 16451 6857
rect 16393 6817 16405 6851
rect 16439 6817 16451 6851
rect 16393 6811 16451 6817
rect 15197 6783 15255 6789
rect 15197 6780 15209 6783
rect 14660 6752 15209 6780
rect 15197 6749 15209 6752
rect 15243 6780 15255 6783
rect 15243 6752 16436 6780
rect 15243 6749 15255 6752
rect 15197 6743 15255 6749
rect 16408 6724 16436 6752
rect 13446 6712 13452 6724
rect 11440 6684 13452 6712
rect 10873 6675 10931 6681
rect 9824 6616 10364 6644
rect 10413 6647 10471 6653
rect 9824 6604 9830 6616
rect 10413 6613 10425 6647
rect 10459 6644 10471 6647
rect 10888 6644 10916 6675
rect 13446 6672 13452 6684
rect 13504 6672 13510 6724
rect 14274 6672 14280 6724
rect 14332 6712 14338 6724
rect 14553 6715 14611 6721
rect 14553 6712 14565 6715
rect 14332 6684 14565 6712
rect 14332 6672 14338 6684
rect 14553 6681 14565 6684
rect 14599 6712 14611 6715
rect 14599 6684 16344 6712
rect 14599 6681 14611 6684
rect 14553 6675 14611 6681
rect 10459 6616 10916 6644
rect 10459 6613 10471 6616
rect 10413 6607 10471 6613
rect 10962 6604 10968 6656
rect 11020 6644 11026 6656
rect 11149 6647 11207 6653
rect 11149 6644 11161 6647
rect 11020 6616 11161 6644
rect 11020 6604 11026 6616
rect 11149 6613 11161 6616
rect 11195 6613 11207 6647
rect 11149 6607 11207 6613
rect 12618 6604 12624 6656
rect 12676 6644 12682 6656
rect 13722 6644 13728 6656
rect 12676 6616 13728 6644
rect 12676 6604 12682 6616
rect 13722 6604 13728 6616
rect 13780 6604 13786 6656
rect 15654 6604 15660 6656
rect 15712 6604 15718 6656
rect 15746 6604 15752 6656
rect 15804 6604 15810 6656
rect 16117 6647 16175 6653
rect 16117 6613 16129 6647
rect 16163 6644 16175 6647
rect 16206 6644 16212 6656
rect 16163 6616 16212 6644
rect 16163 6613 16175 6616
rect 16117 6607 16175 6613
rect 16206 6604 16212 6616
rect 16264 6604 16270 6656
rect 16316 6644 16344 6684
rect 16390 6672 16396 6724
rect 16448 6672 16454 6724
rect 16660 6715 16718 6721
rect 16660 6681 16672 6715
rect 16706 6712 16718 6715
rect 16850 6712 16856 6724
rect 16706 6684 16856 6712
rect 16706 6681 16718 6684
rect 16660 6675 16718 6681
rect 16850 6672 16856 6684
rect 16908 6672 16914 6724
rect 17494 6644 17500 6656
rect 16316 6616 17500 6644
rect 17494 6604 17500 6616
rect 17552 6644 17558 6656
rect 17773 6647 17831 6653
rect 17773 6644 17785 6647
rect 17552 6616 17785 6644
rect 17552 6604 17558 6616
rect 17773 6613 17785 6616
rect 17819 6613 17831 6647
rect 17773 6607 17831 6613
rect 1104 6554 18124 6576
rect 1104 6502 3737 6554
rect 3789 6502 3801 6554
rect 3853 6502 3865 6554
rect 3917 6502 3929 6554
rect 3981 6502 3993 6554
rect 4045 6502 7992 6554
rect 8044 6502 8056 6554
rect 8108 6502 8120 6554
rect 8172 6502 8184 6554
rect 8236 6502 8248 6554
rect 8300 6502 12247 6554
rect 12299 6502 12311 6554
rect 12363 6502 12375 6554
rect 12427 6502 12439 6554
rect 12491 6502 12503 6554
rect 12555 6502 16502 6554
rect 16554 6502 16566 6554
rect 16618 6502 16630 6554
rect 16682 6502 16694 6554
rect 16746 6502 16758 6554
rect 16810 6502 18124 6554
rect 1104 6480 18124 6502
rect 2498 6400 2504 6452
rect 2556 6400 2562 6452
rect 3329 6443 3387 6449
rect 3329 6409 3341 6443
rect 3375 6440 3387 6443
rect 4157 6443 4215 6449
rect 4157 6440 4169 6443
rect 3375 6412 4169 6440
rect 3375 6409 3387 6412
rect 3329 6403 3387 6409
rect 4157 6409 4169 6412
rect 4203 6440 4215 6443
rect 4246 6440 4252 6452
rect 4203 6412 4252 6440
rect 4203 6409 4215 6412
rect 4157 6403 4215 6409
rect 4246 6400 4252 6412
rect 4304 6400 4310 6452
rect 4522 6400 4528 6452
rect 4580 6400 4586 6452
rect 4982 6400 4988 6452
rect 5040 6400 5046 6452
rect 5442 6400 5448 6452
rect 5500 6400 5506 6452
rect 6914 6400 6920 6452
rect 6972 6440 6978 6452
rect 7926 6440 7932 6452
rect 6972 6412 7932 6440
rect 6972 6400 6978 6412
rect 7926 6400 7932 6412
rect 7984 6400 7990 6452
rect 8248 6400 8254 6452
rect 8306 6440 8312 6452
rect 8386 6440 8392 6452
rect 8306 6412 8392 6440
rect 8306 6400 8312 6412
rect 8386 6400 8392 6412
rect 8444 6400 8450 6452
rect 9122 6400 9128 6452
rect 9180 6400 9186 6452
rect 10778 6400 10784 6452
rect 10836 6440 10842 6452
rect 11609 6443 11667 6449
rect 11609 6440 11621 6443
rect 10836 6412 11621 6440
rect 10836 6400 10842 6412
rect 11609 6409 11621 6412
rect 11655 6409 11667 6443
rect 11609 6403 11667 6409
rect 15654 6400 15660 6452
rect 15712 6400 15718 6452
rect 16485 6443 16543 6449
rect 16485 6409 16497 6443
rect 16531 6409 16543 6443
rect 16485 6403 16543 6409
rect 16669 6443 16727 6449
rect 16669 6409 16681 6443
rect 16715 6440 16727 6443
rect 16850 6440 16856 6452
rect 16715 6412 16856 6440
rect 16715 6409 16727 6412
rect 16669 6403 16727 6409
rect 6733 6375 6791 6381
rect 6733 6372 6745 6375
rect 3712 6344 6745 6372
rect 2685 6307 2743 6313
rect 2685 6273 2697 6307
rect 2731 6304 2743 6307
rect 2866 6304 2872 6316
rect 2731 6276 2872 6304
rect 2731 6273 2743 6276
rect 2685 6267 2743 6273
rect 2866 6264 2872 6276
rect 2924 6264 2930 6316
rect 3418 6304 3424 6316
rect 3160 6276 3424 6304
rect 3160 6245 3188 6276
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 3145 6239 3203 6245
rect 3145 6205 3157 6239
rect 3191 6205 3203 6239
rect 3145 6199 3203 6205
rect 3237 6239 3295 6245
rect 3237 6205 3249 6239
rect 3283 6205 3295 6239
rect 3237 6199 3295 6205
rect 3252 6100 3280 6199
rect 3712 6177 3740 6344
rect 6733 6341 6745 6344
rect 6779 6341 6791 6375
rect 6733 6335 6791 6341
rect 7024 6344 8147 6372
rect 4890 6304 4896 6316
rect 3988 6276 4896 6304
rect 3988 6245 4016 6276
rect 4890 6264 4896 6276
rect 4948 6264 4954 6316
rect 6546 6313 6552 6316
rect 5077 6307 5135 6313
rect 5077 6273 5089 6307
rect 5123 6304 5135 6307
rect 5537 6307 5595 6313
rect 5537 6304 5549 6307
rect 5123 6276 5549 6304
rect 5123 6273 5135 6276
rect 5077 6267 5135 6273
rect 5537 6273 5549 6276
rect 5583 6273 5595 6307
rect 6544 6304 6552 6313
rect 6507 6276 6552 6304
rect 5537 6267 5595 6273
rect 6544 6267 6552 6276
rect 6546 6264 6552 6267
rect 6604 6264 6610 6316
rect 6638 6264 6644 6316
rect 6696 6264 6702 6316
rect 6914 6313 6920 6316
rect 6888 6307 6920 6313
rect 6888 6273 6900 6307
rect 6888 6267 6920 6273
rect 6914 6264 6920 6267
rect 6972 6264 6978 6316
rect 7024 6313 7052 6344
rect 7009 6307 7067 6313
rect 7009 6273 7021 6307
rect 7055 6273 7067 6307
rect 7009 6267 7067 6273
rect 7558 6264 7564 6316
rect 7616 6264 7622 6316
rect 7742 6264 7748 6316
rect 7800 6304 7806 6316
rect 8021 6307 8079 6313
rect 8021 6304 8033 6307
rect 7800 6276 8033 6304
rect 7800 6264 7806 6276
rect 8021 6273 8033 6276
rect 8067 6273 8079 6307
rect 8119 6304 8147 6344
rect 8266 6344 10916 6372
rect 8119 6302 8156 6304
rect 8266 6302 8294 6344
rect 8119 6276 8294 6302
rect 8128 6274 8294 6276
rect 8021 6267 8079 6273
rect 8938 6264 8944 6316
rect 8996 6264 9002 6316
rect 10704 6313 10732 6344
rect 10689 6307 10747 6313
rect 10689 6273 10701 6307
rect 10735 6273 10747 6307
rect 10689 6267 10747 6273
rect 10782 6307 10840 6313
rect 10782 6273 10794 6307
rect 10828 6273 10840 6307
rect 10782 6267 10840 6273
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6205 4031 6239
rect 3973 6199 4031 6205
rect 4065 6239 4123 6245
rect 4065 6205 4077 6239
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 3697 6171 3755 6177
rect 3697 6137 3709 6171
rect 3743 6137 3755 6171
rect 3697 6131 3755 6137
rect 4080 6112 4108 6199
rect 4798 6196 4804 6248
rect 4856 6196 4862 6248
rect 6178 6196 6184 6248
rect 6236 6196 6242 6248
rect 7653 6239 7711 6245
rect 7653 6205 7665 6239
rect 7699 6236 7711 6239
rect 7834 6236 7840 6248
rect 7699 6208 7840 6236
rect 7699 6205 7711 6208
rect 7653 6199 7711 6205
rect 7834 6196 7840 6208
rect 7892 6196 7898 6248
rect 7926 6196 7932 6248
rect 7984 6236 7990 6248
rect 10796 6236 10824 6267
rect 7984 6208 10824 6236
rect 7984 6196 7990 6208
rect 6730 6128 6736 6180
rect 6788 6168 6794 6180
rect 7101 6171 7159 6177
rect 7101 6168 7113 6171
rect 6788 6140 7113 6168
rect 6788 6128 6794 6140
rect 7101 6137 7113 6140
rect 7147 6137 7159 6171
rect 7101 6131 7159 6137
rect 7374 6128 7380 6180
rect 7432 6168 7438 6180
rect 9766 6168 9772 6180
rect 7432 6140 9772 6168
rect 7432 6128 7438 6140
rect 9766 6128 9772 6140
rect 9824 6128 9830 6180
rect 10888 6168 10916 6344
rect 11054 6332 11060 6384
rect 11112 6332 11118 6384
rect 12069 6375 12127 6381
rect 12069 6341 12081 6375
rect 12115 6372 12127 6375
rect 13262 6372 13268 6384
rect 12115 6344 13268 6372
rect 12115 6341 12127 6344
rect 12069 6335 12127 6341
rect 13262 6332 13268 6344
rect 13320 6332 13326 6384
rect 15286 6332 15292 6384
rect 15344 6372 15350 6384
rect 15562 6372 15568 6384
rect 15344 6344 15568 6372
rect 15344 6332 15350 6344
rect 15562 6332 15568 6344
rect 15620 6372 15626 6384
rect 16025 6375 16083 6381
rect 16025 6372 16037 6375
rect 15620 6344 16037 6372
rect 15620 6332 15626 6344
rect 16025 6341 16037 6344
rect 16071 6341 16083 6375
rect 16025 6335 16083 6341
rect 10965 6307 11023 6313
rect 10965 6273 10977 6307
rect 11011 6273 11023 6307
rect 10965 6267 11023 6273
rect 10980 6236 11008 6267
rect 11146 6264 11152 6316
rect 11204 6313 11210 6316
rect 11204 6304 11212 6313
rect 11977 6307 12035 6313
rect 11204 6276 11249 6304
rect 11204 6267 11212 6276
rect 11977 6273 11989 6307
rect 12023 6304 12035 6307
rect 12434 6304 12440 6316
rect 12023 6276 12440 6304
rect 12023 6273 12035 6276
rect 11977 6267 12035 6273
rect 11204 6264 11210 6267
rect 12434 6264 12440 6276
rect 12492 6264 12498 6316
rect 12618 6264 12624 6316
rect 12676 6264 12682 6316
rect 15010 6264 15016 6316
rect 15068 6264 15074 6316
rect 16117 6307 16175 6313
rect 16117 6273 16129 6307
rect 16163 6304 16175 6307
rect 16298 6304 16304 6316
rect 16163 6276 16304 6304
rect 16163 6273 16175 6276
rect 16117 6267 16175 6273
rect 16298 6264 16304 6276
rect 16356 6264 16362 6316
rect 16500 6304 16528 6403
rect 16850 6400 16856 6412
rect 16908 6400 16914 6452
rect 16853 6307 16911 6313
rect 16853 6304 16865 6307
rect 16500 6276 16865 6304
rect 16853 6273 16865 6276
rect 16899 6273 16911 6307
rect 16853 6267 16911 6273
rect 17770 6264 17776 6316
rect 17828 6264 17834 6316
rect 11330 6236 11336 6248
rect 10980 6208 11336 6236
rect 11330 6196 11336 6208
rect 11388 6196 11394 6248
rect 12250 6196 12256 6248
rect 12308 6236 12314 6248
rect 14090 6236 14096 6248
rect 12308 6208 14096 6236
rect 12308 6196 12314 6208
rect 14090 6196 14096 6208
rect 14148 6196 14154 6248
rect 15470 6196 15476 6248
rect 15528 6236 15534 6248
rect 15838 6236 15844 6248
rect 15528 6208 15844 6236
rect 15528 6196 15534 6208
rect 15838 6196 15844 6208
rect 15896 6196 15902 6248
rect 16390 6196 16396 6248
rect 16448 6236 16454 6248
rect 17497 6239 17555 6245
rect 17497 6236 17509 6239
rect 16448 6208 17509 6236
rect 16448 6196 16454 6208
rect 17497 6205 17509 6208
rect 17543 6205 17555 6239
rect 17497 6199 17555 6205
rect 13078 6168 13084 6180
rect 10888 6140 13084 6168
rect 13078 6128 13084 6140
rect 13136 6128 13142 6180
rect 4062 6100 4068 6112
rect 3252 6072 4068 6100
rect 4062 6060 4068 6072
rect 4120 6060 4126 6112
rect 6270 6060 6276 6112
rect 6328 6100 6334 6112
rect 6365 6103 6423 6109
rect 6365 6100 6377 6103
rect 6328 6072 6377 6100
rect 6328 6060 6334 6072
rect 6365 6069 6377 6072
rect 6411 6069 6423 6103
rect 6365 6063 6423 6069
rect 7282 6060 7288 6112
rect 7340 6060 7346 6112
rect 8110 6060 8116 6112
rect 8168 6100 8174 6112
rect 8205 6103 8263 6109
rect 8205 6100 8217 6103
rect 8168 6072 8217 6100
rect 8168 6060 8174 6072
rect 8205 6069 8217 6072
rect 8251 6069 8263 6103
rect 8205 6063 8263 6069
rect 11333 6103 11391 6109
rect 11333 6069 11345 6103
rect 11379 6100 11391 6103
rect 11422 6100 11428 6112
rect 11379 6072 11428 6100
rect 11379 6069 11391 6072
rect 11333 6063 11391 6069
rect 11422 6060 11428 6072
rect 11480 6060 11486 6112
rect 1104 6010 18124 6032
rect 1104 5958 3077 6010
rect 3129 5958 3141 6010
rect 3193 5958 3205 6010
rect 3257 5958 3269 6010
rect 3321 5958 3333 6010
rect 3385 5958 7332 6010
rect 7384 5958 7396 6010
rect 7448 5958 7460 6010
rect 7512 5958 7524 6010
rect 7576 5958 7588 6010
rect 7640 5958 11587 6010
rect 11639 5958 11651 6010
rect 11703 5958 11715 6010
rect 11767 5958 11779 6010
rect 11831 5958 11843 6010
rect 11895 5958 15842 6010
rect 15894 5958 15906 6010
rect 15958 5958 15970 6010
rect 16022 5958 16034 6010
rect 16086 5958 16098 6010
rect 16150 5958 18124 6010
rect 1104 5936 18124 5958
rect 3605 5899 3663 5905
rect 3605 5865 3617 5899
rect 3651 5896 3663 5899
rect 4338 5896 4344 5908
rect 3651 5868 4344 5896
rect 3651 5865 3663 5868
rect 3605 5859 3663 5865
rect 4338 5856 4344 5868
rect 4396 5856 4402 5908
rect 5813 5899 5871 5905
rect 5813 5865 5825 5899
rect 5859 5865 5871 5899
rect 5813 5859 5871 5865
rect 5997 5899 6055 5905
rect 5997 5865 6009 5899
rect 6043 5896 6055 5899
rect 6638 5896 6644 5908
rect 6043 5868 6644 5896
rect 6043 5865 6055 5868
rect 5997 5859 6055 5865
rect 3418 5788 3424 5840
rect 3476 5828 3482 5840
rect 3789 5831 3847 5837
rect 3789 5828 3801 5831
rect 3476 5800 3801 5828
rect 3476 5788 3482 5800
rect 3789 5797 3801 5800
rect 3835 5797 3847 5831
rect 3789 5791 3847 5797
rect 4062 5788 4068 5840
rect 4120 5828 4126 5840
rect 5828 5828 5856 5859
rect 6638 5856 6644 5868
rect 6696 5856 6702 5908
rect 7392 5868 10732 5896
rect 6178 5828 6184 5840
rect 4120 5800 5212 5828
rect 5828 5800 6184 5828
rect 4120 5788 4126 5800
rect 4430 5720 4436 5772
rect 4488 5720 4494 5772
rect 5184 5769 5212 5800
rect 6178 5788 6184 5800
rect 6236 5788 6242 5840
rect 7006 5788 7012 5840
rect 7064 5828 7070 5840
rect 7064 5800 7144 5828
rect 7064 5788 7070 5800
rect 5169 5763 5227 5769
rect 5169 5729 5181 5763
rect 5215 5729 5227 5763
rect 5169 5723 5227 5729
rect 6549 5763 6607 5769
rect 6549 5729 6561 5763
rect 6595 5760 6607 5763
rect 6914 5760 6920 5772
rect 6595 5732 6920 5760
rect 6595 5729 6607 5732
rect 6549 5723 6607 5729
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 7116 5769 7144 5800
rect 7101 5763 7159 5769
rect 7101 5729 7113 5763
rect 7147 5760 7159 5763
rect 7392 5760 7420 5868
rect 8757 5831 8815 5837
rect 8757 5797 8769 5831
rect 8803 5828 8815 5831
rect 10704 5828 10732 5868
rect 11330 5856 11336 5908
rect 11388 5896 11394 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 11388 5868 12817 5896
rect 11388 5856 11394 5868
rect 12805 5865 12817 5868
rect 12851 5865 12863 5899
rect 12805 5859 12863 5865
rect 14918 5856 14924 5908
rect 14976 5856 14982 5908
rect 13446 5828 13452 5840
rect 8803 5800 9536 5828
rect 8803 5797 8815 5800
rect 8757 5791 8815 5797
rect 9508 5772 9536 5800
rect 10704 5800 13452 5828
rect 7147 5732 7420 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 9490 5720 9496 5772
rect 9548 5720 9554 5772
rect 10704 5769 10732 5800
rect 13446 5788 13452 5800
rect 13504 5788 13510 5840
rect 15378 5788 15384 5840
rect 15436 5828 15442 5840
rect 16393 5831 16451 5837
rect 15436 5800 15792 5828
rect 15436 5788 15442 5800
rect 10689 5763 10747 5769
rect 10689 5729 10701 5763
rect 10735 5729 10747 5763
rect 10689 5723 10747 5729
rect 10781 5763 10839 5769
rect 10781 5729 10793 5763
rect 10827 5760 10839 5763
rect 11054 5760 11060 5772
rect 10827 5732 11060 5760
rect 10827 5729 10839 5732
rect 10781 5723 10839 5729
rect 11054 5720 11060 5732
rect 11112 5720 11118 5772
rect 11146 5720 11152 5772
rect 11204 5760 11210 5772
rect 11333 5763 11391 5769
rect 11333 5760 11345 5763
rect 11204 5732 11345 5760
rect 11204 5720 11210 5732
rect 11333 5729 11345 5732
rect 11379 5729 11391 5763
rect 12986 5760 12992 5772
rect 11333 5723 11391 5729
rect 11808 5732 12992 5760
rect 3421 5695 3479 5701
rect 3421 5661 3433 5695
rect 3467 5692 3479 5695
rect 4522 5692 4528 5704
rect 3467 5664 4528 5692
rect 3467 5661 3479 5664
rect 3421 5655 3479 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 5534 5652 5540 5704
rect 5592 5652 5598 5704
rect 6270 5652 6276 5704
rect 6328 5652 6334 5704
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 6822 5652 6828 5704
rect 6880 5652 6886 5704
rect 7006 5652 7012 5704
rect 7064 5652 7070 5704
rect 7377 5695 7435 5701
rect 7377 5661 7389 5695
rect 7423 5692 7435 5695
rect 7423 5664 7880 5692
rect 7423 5661 7435 5664
rect 7377 5655 7435 5661
rect 7852 5636 7880 5664
rect 10962 5652 10968 5704
rect 11020 5652 11026 5704
rect 11238 5652 11244 5704
rect 11296 5652 11302 5704
rect 11422 5652 11428 5704
rect 11480 5692 11486 5704
rect 11517 5695 11575 5701
rect 11517 5692 11529 5695
rect 11480 5664 11529 5692
rect 11480 5652 11486 5664
rect 11517 5661 11529 5664
rect 11563 5661 11575 5695
rect 11517 5655 11575 5661
rect 4157 5627 4215 5633
rect 4157 5593 4169 5627
rect 4203 5624 4215 5627
rect 4617 5627 4675 5633
rect 4617 5624 4629 5627
rect 4203 5596 4629 5624
rect 4203 5593 4215 5596
rect 4157 5587 4215 5593
rect 4617 5593 4629 5596
rect 4663 5593 4675 5627
rect 4617 5587 4675 5593
rect 7644 5627 7702 5633
rect 7644 5593 7656 5627
rect 7690 5624 7702 5627
rect 7742 5624 7748 5636
rect 7690 5596 7748 5624
rect 7690 5593 7702 5596
rect 7644 5587 7702 5593
rect 7742 5584 7748 5596
rect 7800 5584 7806 5636
rect 7834 5584 7840 5636
rect 7892 5584 7898 5636
rect 11149 5627 11207 5633
rect 11149 5593 11161 5627
rect 11195 5624 11207 5627
rect 11808 5624 11836 5732
rect 12986 5720 12992 5732
rect 13044 5720 13050 5772
rect 13262 5720 13268 5772
rect 13320 5720 13326 5772
rect 13357 5763 13415 5769
rect 13357 5729 13369 5763
rect 13403 5760 13415 5763
rect 13538 5760 13544 5772
rect 13403 5732 13544 5760
rect 13403 5729 13415 5732
rect 13357 5723 13415 5729
rect 13538 5720 13544 5732
rect 13596 5720 13602 5772
rect 14366 5720 14372 5772
rect 14424 5720 14430 5772
rect 15654 5760 15660 5772
rect 14476 5732 15660 5760
rect 12250 5652 12256 5704
rect 12308 5652 12314 5704
rect 12434 5652 12440 5704
rect 12492 5692 12498 5704
rect 13173 5695 13231 5701
rect 13173 5692 13185 5695
rect 12492 5664 13185 5692
rect 12492 5652 12498 5664
rect 13173 5661 13185 5664
rect 13219 5692 13231 5695
rect 14476 5692 14504 5732
rect 15654 5720 15660 5732
rect 15712 5720 15718 5772
rect 15764 5769 15792 5800
rect 16393 5797 16405 5831
rect 16439 5797 16451 5831
rect 16393 5791 16451 5797
rect 15749 5763 15807 5769
rect 15749 5729 15761 5763
rect 15795 5729 15807 5763
rect 15749 5723 15807 5729
rect 15838 5720 15844 5772
rect 15896 5760 15902 5772
rect 15933 5763 15991 5769
rect 15933 5760 15945 5763
rect 15896 5732 15945 5760
rect 15896 5720 15902 5732
rect 15933 5729 15945 5732
rect 15979 5729 15991 5763
rect 15933 5723 15991 5729
rect 13219 5664 14504 5692
rect 13219 5661 13231 5664
rect 13173 5655 13231 5661
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 15378 5652 15384 5704
rect 15436 5652 15442 5704
rect 16408 5692 16436 5791
rect 17770 5720 17776 5772
rect 17828 5720 17834 5772
rect 16485 5695 16543 5701
rect 16485 5692 16497 5695
rect 16408 5664 16497 5692
rect 16485 5661 16497 5664
rect 16531 5661 16543 5695
rect 16485 5655 16543 5661
rect 17497 5695 17555 5701
rect 17497 5661 17509 5695
rect 17543 5661 17555 5695
rect 17497 5655 17555 5661
rect 11195 5596 11836 5624
rect 12529 5627 12587 5633
rect 11195 5593 11207 5596
rect 11149 5587 11207 5593
rect 12529 5593 12541 5627
rect 12575 5624 12587 5627
rect 12710 5624 12716 5636
rect 12575 5596 12716 5624
rect 12575 5593 12587 5596
rect 12529 5587 12587 5593
rect 12710 5584 12716 5596
rect 12768 5584 12774 5636
rect 13538 5584 13544 5636
rect 13596 5624 13602 5636
rect 14568 5624 14596 5652
rect 15013 5627 15071 5633
rect 15013 5624 15025 5627
rect 13596 5596 15025 5624
rect 13596 5584 13602 5596
rect 15013 5593 15025 5596
rect 15059 5624 15071 5627
rect 15059 5596 15332 5624
rect 15059 5593 15071 5596
rect 15013 5587 15071 5593
rect 4249 5559 4307 5565
rect 4249 5525 4261 5559
rect 4295 5556 4307 5559
rect 4982 5556 4988 5568
rect 4295 5528 4988 5556
rect 4295 5525 4307 5528
rect 4249 5519 4307 5525
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 6086 5516 6092 5568
rect 6144 5516 6150 5568
rect 6270 5516 6276 5568
rect 6328 5556 6334 5568
rect 6641 5559 6699 5565
rect 6641 5556 6653 5559
rect 6328 5528 6653 5556
rect 6328 5516 6334 5528
rect 6641 5525 6653 5528
rect 6687 5525 6699 5559
rect 6641 5519 6699 5525
rect 8938 5516 8944 5568
rect 8996 5516 9002 5568
rect 11701 5559 11759 5565
rect 11701 5525 11713 5559
rect 11747 5556 11759 5559
rect 13354 5556 13360 5568
rect 11747 5528 13360 5556
rect 11747 5525 11759 5528
rect 11701 5519 11759 5525
rect 13354 5516 13360 5528
rect 13412 5516 13418 5568
rect 15194 5516 15200 5568
rect 15252 5516 15258 5568
rect 15304 5556 15332 5596
rect 15746 5584 15752 5636
rect 15804 5624 15810 5636
rect 16025 5627 16083 5633
rect 16025 5624 16037 5627
rect 15804 5596 16037 5624
rect 15804 5584 15810 5596
rect 16025 5593 16037 5596
rect 16071 5593 16083 5627
rect 17512 5624 17540 5655
rect 16025 5587 16083 5593
rect 16132 5596 17540 5624
rect 16132 5556 16160 5596
rect 15304 5528 16160 5556
rect 16669 5559 16727 5565
rect 16669 5525 16681 5559
rect 16715 5556 16727 5559
rect 17034 5556 17040 5568
rect 16715 5528 17040 5556
rect 16715 5525 16727 5528
rect 16669 5519 16727 5525
rect 17034 5516 17040 5528
rect 17092 5516 17098 5568
rect 1104 5466 18124 5488
rect 1104 5414 3737 5466
rect 3789 5414 3801 5466
rect 3853 5414 3865 5466
rect 3917 5414 3929 5466
rect 3981 5414 3993 5466
rect 4045 5414 7992 5466
rect 8044 5414 8056 5466
rect 8108 5414 8120 5466
rect 8172 5414 8184 5466
rect 8236 5414 8248 5466
rect 8300 5414 12247 5466
rect 12299 5414 12311 5466
rect 12363 5414 12375 5466
rect 12427 5414 12439 5466
rect 12491 5414 12503 5466
rect 12555 5414 16502 5466
rect 16554 5414 16566 5466
rect 16618 5414 16630 5466
rect 16682 5414 16694 5466
rect 16746 5414 16758 5466
rect 16810 5414 18124 5466
rect 1104 5392 18124 5414
rect 3973 5355 4031 5361
rect 3973 5321 3985 5355
rect 4019 5352 4031 5355
rect 4062 5352 4068 5364
rect 4019 5324 4068 5352
rect 4019 5321 4031 5324
rect 3973 5315 4031 5321
rect 4062 5312 4068 5324
rect 4120 5312 4126 5364
rect 7006 5312 7012 5364
rect 7064 5352 7070 5364
rect 8205 5355 8263 5361
rect 8205 5352 8217 5355
rect 7064 5324 8217 5352
rect 7064 5312 7070 5324
rect 8205 5321 8217 5324
rect 8251 5321 8263 5355
rect 8205 5315 8263 5321
rect 8757 5355 8815 5361
rect 8757 5321 8769 5355
rect 8803 5352 8815 5355
rect 8938 5352 8944 5364
rect 8803 5324 8944 5352
rect 8803 5321 8815 5324
rect 8757 5315 8815 5321
rect 8938 5312 8944 5324
rect 8996 5312 9002 5364
rect 9030 5312 9036 5364
rect 9088 5352 9094 5364
rect 10410 5352 10416 5364
rect 9088 5324 10416 5352
rect 9088 5312 9094 5324
rect 10410 5312 10416 5324
rect 10468 5352 10474 5364
rect 10962 5352 10968 5364
rect 10468 5324 10968 5352
rect 10468 5312 10474 5324
rect 10962 5312 10968 5324
rect 11020 5312 11026 5364
rect 11054 5312 11060 5364
rect 11112 5312 11118 5364
rect 13262 5312 13268 5364
rect 13320 5352 13326 5364
rect 16117 5355 16175 5361
rect 16117 5352 16129 5355
rect 13320 5324 16129 5352
rect 13320 5312 13326 5324
rect 16117 5321 16129 5324
rect 16163 5321 16175 5355
rect 16117 5315 16175 5321
rect 4338 5293 4344 5296
rect 4332 5284 4344 5293
rect 2608 5256 4108 5284
rect 4299 5256 4344 5284
rect 2608 5225 2636 5256
rect 2866 5225 2872 5228
rect 2593 5219 2651 5225
rect 2593 5185 2605 5219
rect 2639 5185 2651 5219
rect 2593 5179 2651 5185
rect 2860 5179 2872 5225
rect 2866 5176 2872 5179
rect 2924 5176 2930 5228
rect 4080 5160 4108 5256
rect 4332 5247 4344 5256
rect 4338 5244 4344 5247
rect 4396 5244 4402 5296
rect 15004 5287 15062 5293
rect 15004 5253 15016 5287
rect 15050 5284 15062 5287
rect 15194 5284 15200 5296
rect 15050 5256 15200 5284
rect 15050 5253 15062 5256
rect 15004 5247 15062 5253
rect 15194 5244 15200 5256
rect 15252 5244 15258 5296
rect 16132 5284 16160 5315
rect 16132 5256 17540 5284
rect 6181 5219 6239 5225
rect 6181 5216 6193 5219
rect 5460 5188 6193 5216
rect 4062 5108 4068 5160
rect 4120 5108 4126 5160
rect 5460 5089 5488 5188
rect 6181 5185 6193 5188
rect 6227 5216 6239 5219
rect 6227 5188 6684 5216
rect 6227 5185 6239 5188
rect 6181 5179 6239 5185
rect 6656 5160 6684 5188
rect 7282 5176 7288 5228
rect 7340 5176 7346 5228
rect 7558 5176 7564 5228
rect 7616 5176 7622 5228
rect 9582 5216 9588 5228
rect 8864 5188 9588 5216
rect 8864 5160 8892 5188
rect 9582 5176 9588 5188
rect 9640 5176 9646 5228
rect 11422 5176 11428 5228
rect 11480 5216 11486 5228
rect 11701 5219 11759 5225
rect 11701 5216 11713 5219
rect 11480 5188 11713 5216
rect 11480 5176 11486 5188
rect 11701 5185 11713 5188
rect 11747 5185 11759 5219
rect 13170 5216 13176 5228
rect 11701 5179 11759 5185
rect 11992 5188 13176 5216
rect 6365 5151 6423 5157
rect 6365 5117 6377 5151
rect 6411 5117 6423 5151
rect 6365 5111 6423 5117
rect 6549 5151 6607 5157
rect 6549 5117 6561 5151
rect 6595 5117 6607 5151
rect 6549 5111 6607 5117
rect 5445 5083 5503 5089
rect 5445 5049 5457 5083
rect 5491 5049 5503 5083
rect 5445 5043 5503 5049
rect 5534 4972 5540 5024
rect 5592 4972 5598 5024
rect 6380 5012 6408 5111
rect 6564 5080 6592 5111
rect 6638 5108 6644 5160
rect 6696 5148 6702 5160
rect 7402 5151 7460 5157
rect 7402 5148 7414 5151
rect 6696 5120 7414 5148
rect 6696 5108 6702 5120
rect 7402 5117 7414 5120
rect 7448 5117 7460 5151
rect 7402 5111 7460 5117
rect 8846 5108 8852 5160
rect 8904 5108 8910 5160
rect 9030 5108 9036 5160
rect 9088 5108 9094 5160
rect 9217 5151 9275 5157
rect 9217 5117 9229 5151
rect 9263 5117 9275 5151
rect 9217 5111 9275 5117
rect 9401 5151 9459 5157
rect 9401 5117 9413 5151
rect 9447 5148 9459 5151
rect 9766 5148 9772 5160
rect 9447 5120 9772 5148
rect 9447 5117 9459 5120
rect 9401 5111 9459 5117
rect 6822 5080 6828 5092
rect 6564 5052 6828 5080
rect 6822 5040 6828 5052
rect 6880 5040 6886 5092
rect 7006 5040 7012 5092
rect 7064 5040 7070 5092
rect 8018 5040 8024 5092
rect 8076 5080 8082 5092
rect 9232 5080 9260 5111
rect 9766 5108 9772 5120
rect 9824 5108 9830 5160
rect 10134 5108 10140 5160
rect 10192 5108 10198 5160
rect 10226 5108 10232 5160
rect 10284 5157 10290 5160
rect 10284 5151 10312 5157
rect 10300 5117 10312 5151
rect 10284 5111 10312 5117
rect 10284 5108 10290 5111
rect 10410 5108 10416 5160
rect 10468 5148 10474 5160
rect 11992 5148 12020 5188
rect 13170 5176 13176 5188
rect 13228 5176 13234 5228
rect 13722 5176 13728 5228
rect 13780 5176 13786 5228
rect 13814 5176 13820 5228
rect 13872 5225 13878 5228
rect 13872 5219 13900 5225
rect 13888 5185 13900 5219
rect 13872 5179 13900 5185
rect 13872 5176 13878 5179
rect 14826 5176 14832 5228
rect 14884 5216 14890 5228
rect 17405 5219 17463 5225
rect 17405 5216 17417 5219
rect 14884 5188 17417 5216
rect 14884 5176 14890 5188
rect 17405 5185 17417 5188
rect 17451 5185 17463 5219
rect 17405 5179 17463 5185
rect 10468 5120 12020 5148
rect 10468 5108 10474 5120
rect 12802 5108 12808 5160
rect 12860 5108 12866 5160
rect 12989 5151 13047 5157
rect 12989 5117 13001 5151
rect 13035 5148 13047 5151
rect 13078 5148 13084 5160
rect 13035 5120 13084 5148
rect 13035 5117 13047 5120
rect 12989 5111 13047 5117
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13188 5148 13216 5176
rect 14001 5151 14059 5157
rect 14001 5148 14013 5151
rect 13188 5120 14013 5148
rect 14001 5117 14013 5120
rect 14047 5117 14059 5151
rect 14001 5111 14059 5117
rect 14642 5108 14648 5160
rect 14700 5148 14706 5160
rect 14737 5151 14795 5157
rect 14737 5148 14749 5151
rect 14700 5120 14749 5148
rect 14700 5108 14706 5120
rect 14737 5117 14749 5120
rect 14783 5117 14795 5151
rect 14737 5111 14795 5117
rect 17313 5151 17371 5157
rect 17313 5117 17325 5151
rect 17359 5148 17371 5151
rect 17512 5148 17540 5256
rect 17359 5120 17540 5148
rect 17359 5117 17371 5120
rect 17313 5111 17371 5117
rect 9674 5080 9680 5092
rect 8076 5052 8524 5080
rect 9232 5052 9680 5080
rect 8076 5040 8082 5052
rect 6914 5012 6920 5024
rect 6380 4984 6920 5012
rect 6914 4972 6920 4984
rect 6972 4972 6978 5024
rect 8294 4972 8300 5024
rect 8352 5012 8358 5024
rect 8389 5015 8447 5021
rect 8389 5012 8401 5015
rect 8352 4984 8401 5012
rect 8352 4972 8358 4984
rect 8389 4981 8401 4984
rect 8435 4981 8447 5015
rect 8496 5012 8524 5052
rect 9674 5040 9680 5052
rect 9732 5040 9738 5092
rect 9861 5083 9919 5089
rect 9861 5049 9873 5083
rect 9907 5049 9919 5083
rect 12710 5080 12716 5092
rect 9861 5043 9919 5049
rect 10796 5052 12716 5080
rect 9876 5012 9904 5043
rect 10796 5012 10824 5052
rect 12710 5040 12716 5052
rect 12768 5080 12774 5092
rect 13449 5083 13507 5089
rect 13449 5080 13461 5083
rect 12768 5052 13461 5080
rect 12768 5040 12774 5052
rect 13449 5049 13461 5052
rect 13495 5049 13507 5083
rect 13449 5043 13507 5049
rect 8496 4984 10824 5012
rect 8389 4975 8447 4981
rect 11330 4972 11336 5024
rect 11388 5012 11394 5024
rect 11517 5015 11575 5021
rect 11517 5012 11529 5015
rect 11388 4984 11529 5012
rect 11388 4972 11394 4984
rect 11517 4981 11529 4984
rect 11563 4981 11575 5015
rect 11517 4975 11575 4981
rect 13538 4972 13544 5024
rect 13596 5012 13602 5024
rect 14645 5015 14703 5021
rect 14645 5012 14657 5015
rect 13596 4984 14657 5012
rect 13596 4972 13602 4984
rect 14645 4981 14657 4984
rect 14691 4981 14703 5015
rect 14645 4975 14703 4981
rect 16206 4972 16212 5024
rect 16264 5012 16270 5024
rect 16669 5015 16727 5021
rect 16669 5012 16681 5015
rect 16264 4984 16681 5012
rect 16264 4972 16270 4984
rect 16669 4981 16681 4984
rect 16715 4981 16727 5015
rect 16669 4975 16727 4981
rect 17586 4972 17592 5024
rect 17644 4972 17650 5024
rect 1104 4922 18124 4944
rect 1104 4870 3077 4922
rect 3129 4870 3141 4922
rect 3193 4870 3205 4922
rect 3257 4870 3269 4922
rect 3321 4870 3333 4922
rect 3385 4870 7332 4922
rect 7384 4870 7396 4922
rect 7448 4870 7460 4922
rect 7512 4870 7524 4922
rect 7576 4870 7588 4922
rect 7640 4870 11587 4922
rect 11639 4870 11651 4922
rect 11703 4870 11715 4922
rect 11767 4870 11779 4922
rect 11831 4870 11843 4922
rect 11895 4870 15842 4922
rect 15894 4870 15906 4922
rect 15958 4870 15970 4922
rect 16022 4870 16034 4922
rect 16086 4870 16098 4922
rect 16150 4870 18124 4922
rect 1104 4848 18124 4870
rect 2866 4768 2872 4820
rect 2924 4808 2930 4820
rect 2961 4811 3019 4817
rect 2961 4808 2973 4811
rect 2924 4780 2973 4808
rect 2924 4768 2930 4780
rect 2961 4777 2973 4780
rect 3007 4777 3019 4811
rect 2961 4771 3019 4777
rect 4522 4768 4528 4820
rect 4580 4768 4586 4820
rect 5629 4811 5687 4817
rect 5629 4777 5641 4811
rect 5675 4808 5687 4811
rect 6454 4808 6460 4820
rect 5675 4780 6460 4808
rect 5675 4777 5687 4780
rect 5629 4771 5687 4777
rect 6454 4768 6460 4780
rect 6512 4768 6518 4820
rect 6546 4768 6552 4820
rect 6604 4808 6610 4820
rect 6604 4780 6868 4808
rect 6604 4768 6610 4780
rect 6840 4749 6868 4780
rect 7006 4768 7012 4820
rect 7064 4808 7070 4820
rect 7064 4780 7420 4808
rect 7064 4768 7070 4780
rect 6825 4743 6883 4749
rect 6825 4709 6837 4743
rect 6871 4709 6883 4743
rect 6825 4703 6883 4709
rect 4982 4632 4988 4684
rect 5040 4632 5046 4684
rect 5166 4632 5172 4684
rect 5224 4632 5230 4684
rect 5902 4632 5908 4684
rect 5960 4672 5966 4684
rect 6263 4675 6321 4681
rect 6263 4672 6275 4675
rect 5960 4644 6275 4672
rect 5960 4632 5966 4644
rect 6263 4641 6275 4644
rect 6309 4641 6321 4675
rect 6263 4635 6321 4641
rect 6530 4675 6588 4681
rect 6530 4641 6542 4675
rect 6576 4672 6588 4675
rect 6730 4672 6736 4684
rect 6576 4644 6736 4672
rect 6576 4641 6588 4644
rect 6530 4635 6588 4641
rect 6730 4632 6736 4644
rect 6788 4632 6794 4684
rect 7392 4672 7420 4780
rect 7742 4768 7748 4820
rect 7800 4808 7806 4820
rect 8113 4811 8171 4817
rect 8113 4808 8125 4811
rect 7800 4780 8125 4808
rect 7800 4768 7806 4780
rect 8113 4777 8125 4780
rect 8159 4777 8171 4811
rect 10410 4808 10416 4820
rect 8113 4771 8171 4777
rect 9416 4780 10416 4808
rect 7650 4700 7656 4752
rect 7708 4740 7714 4752
rect 9416 4740 9444 4780
rect 10410 4768 10416 4780
rect 10468 4768 10474 4820
rect 11057 4811 11115 4817
rect 11057 4777 11069 4811
rect 11103 4808 11115 4811
rect 11146 4808 11152 4820
rect 11103 4780 11152 4808
rect 11103 4777 11115 4780
rect 11057 4771 11115 4777
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 13538 4768 13544 4820
rect 13596 4768 13602 4820
rect 13909 4811 13967 4817
rect 13909 4777 13921 4811
rect 13955 4808 13967 4811
rect 14826 4808 14832 4820
rect 13955 4780 14832 4808
rect 13955 4777 13967 4780
rect 13909 4771 13967 4777
rect 14826 4768 14832 4780
rect 14884 4768 14890 4820
rect 15013 4811 15071 4817
rect 15013 4777 15025 4811
rect 15059 4808 15071 4811
rect 15378 4808 15384 4820
rect 15059 4780 15384 4808
rect 15059 4777 15071 4780
rect 15013 4771 15071 4777
rect 15378 4768 15384 4780
rect 15436 4768 15442 4820
rect 15488 4780 17540 4808
rect 7708 4712 9444 4740
rect 7708 4700 7714 4712
rect 9490 4700 9496 4752
rect 9548 4740 9554 4752
rect 12621 4743 12679 4749
rect 9548 4712 9996 4740
rect 9548 4700 9554 4712
rect 7469 4675 7527 4681
rect 7469 4672 7481 4675
rect 7392 4644 7481 4672
rect 7469 4641 7481 4644
rect 7515 4672 7527 4675
rect 7742 4672 7748 4684
rect 7515 4644 7748 4672
rect 7515 4641 7527 4644
rect 7469 4635 7527 4641
rect 7742 4632 7748 4644
rect 7800 4632 7806 4684
rect 9401 4675 9459 4681
rect 9401 4641 9413 4675
rect 9447 4672 9459 4675
rect 9766 4672 9772 4684
rect 9447 4644 9772 4672
rect 9447 4641 9459 4644
rect 9401 4635 9459 4641
rect 9766 4632 9772 4644
rect 9824 4632 9830 4684
rect 9858 4632 9864 4684
rect 9916 4632 9922 4684
rect 9968 4672 9996 4712
rect 12621 4709 12633 4743
rect 12667 4709 12679 4743
rect 12621 4703 12679 4709
rect 14921 4743 14979 4749
rect 14921 4709 14933 4743
rect 14967 4740 14979 4743
rect 15488 4740 15516 4780
rect 16206 4740 16212 4752
rect 14967 4712 15516 4740
rect 15580 4712 16212 4740
rect 14967 4709 14979 4712
rect 14921 4703 14979 4709
rect 10226 4672 10232 4684
rect 10284 4681 10290 4684
rect 10284 4675 10312 4681
rect 9968 4644 10232 4672
rect 10226 4632 10232 4644
rect 10300 4641 10312 4675
rect 10284 4635 10312 4641
rect 10284 4632 10290 4635
rect 10410 4632 10416 4684
rect 10468 4672 10474 4684
rect 12636 4672 12664 4703
rect 13357 4675 13415 4681
rect 13357 4672 13369 4675
rect 10468 4644 11008 4672
rect 12636 4644 13369 4672
rect 10468 4632 10474 4644
rect 3145 4607 3203 4613
rect 3145 4573 3157 4607
rect 3191 4604 3203 4607
rect 3418 4604 3424 4616
rect 3191 4576 3424 4604
rect 3191 4573 3203 4576
rect 3145 4567 3203 4573
rect 3418 4564 3424 4576
rect 3476 4564 3482 4616
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 5534 4604 5540 4616
rect 4939 4576 5540 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 5534 4564 5540 4576
rect 5592 4564 5598 4616
rect 6362 4564 6368 4616
rect 6420 4613 6426 4616
rect 6420 4607 6469 4613
rect 6420 4573 6423 4607
rect 6457 4573 6469 4607
rect 6420 4567 6469 4573
rect 6420 4564 6426 4567
rect 7282 4564 7288 4616
rect 7340 4564 7346 4616
rect 8294 4564 8300 4616
rect 8352 4564 8358 4616
rect 9217 4607 9275 4613
rect 9217 4573 9229 4607
rect 9263 4604 9275 4607
rect 9263 4576 9444 4604
rect 9263 4573 9275 4576
rect 9217 4567 9275 4573
rect 6914 4428 6920 4480
rect 6972 4468 6978 4480
rect 7374 4468 7380 4480
rect 6972 4440 7380 4468
rect 6972 4428 6978 4440
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 9416 4468 9444 4576
rect 10134 4564 10140 4616
rect 10192 4564 10198 4616
rect 9674 4468 9680 4480
rect 9416 4440 9680 4468
rect 9674 4428 9680 4440
rect 9732 4468 9738 4480
rect 10410 4468 10416 4480
rect 9732 4440 10416 4468
rect 9732 4428 9738 4440
rect 10410 4428 10416 4440
rect 10468 4428 10474 4480
rect 10980 4468 11008 4644
rect 13357 4641 13369 4644
rect 13403 4672 13415 4675
rect 13814 4672 13820 4684
rect 13403 4644 13820 4672
rect 13403 4641 13415 4644
rect 13357 4635 13415 4641
rect 13814 4632 13820 4644
rect 13872 4632 13878 4684
rect 14182 4632 14188 4684
rect 14240 4672 14246 4684
rect 14240 4644 14780 4672
rect 14240 4632 14246 4644
rect 11241 4607 11299 4613
rect 11241 4573 11253 4607
rect 11287 4604 11299 4607
rect 12618 4604 12624 4616
rect 11287 4576 12624 4604
rect 11287 4573 11299 4576
rect 11241 4567 11299 4573
rect 12618 4564 12624 4576
rect 12676 4564 12682 4616
rect 13446 4564 13452 4616
rect 13504 4564 13510 4616
rect 13630 4564 13636 4616
rect 13688 4604 13694 4616
rect 13725 4607 13783 4613
rect 13725 4604 13737 4607
rect 13688 4576 13737 4604
rect 13688 4564 13694 4576
rect 13725 4573 13737 4576
rect 13771 4573 13783 4607
rect 13725 4567 13783 4573
rect 14458 4564 14464 4616
rect 14516 4564 14522 4616
rect 14550 4564 14556 4616
rect 14608 4564 14614 4616
rect 14752 4613 14780 4644
rect 14737 4607 14795 4613
rect 14737 4573 14749 4607
rect 14783 4573 14795 4607
rect 14737 4567 14795 4573
rect 15381 4607 15439 4613
rect 15381 4573 15393 4607
rect 15427 4604 15439 4607
rect 15580 4604 15608 4712
rect 16206 4700 16212 4712
rect 16264 4700 16270 4752
rect 15657 4675 15715 4681
rect 15657 4641 15669 4675
rect 15703 4672 15715 4675
rect 15838 4672 15844 4684
rect 15703 4644 15844 4672
rect 15703 4641 15715 4644
rect 15657 4635 15715 4641
rect 15838 4632 15844 4644
rect 15896 4632 15902 4684
rect 17512 4613 17540 4780
rect 17678 4768 17684 4820
rect 17736 4768 17742 4820
rect 17313 4607 17371 4613
rect 17313 4604 17325 4607
rect 15427 4576 15608 4604
rect 15672 4576 17325 4604
rect 15427 4573 15439 4576
rect 15381 4567 15439 4573
rect 11330 4496 11336 4548
rect 11388 4536 11394 4548
rect 11486 4539 11544 4545
rect 11486 4536 11498 4539
rect 11388 4508 11498 4536
rect 11388 4496 11394 4508
rect 11486 4505 11498 4508
rect 11532 4505 11544 4539
rect 13998 4536 14004 4548
rect 11486 4499 11544 4505
rect 12406 4508 14004 4536
rect 12406 4468 12434 4508
rect 13998 4496 14004 4508
rect 14056 4496 14062 4548
rect 14642 4496 14648 4548
rect 14700 4536 14706 4548
rect 15672 4536 15700 4576
rect 17313 4573 17325 4576
rect 17359 4573 17371 4607
rect 17313 4567 17371 4573
rect 17497 4607 17555 4613
rect 17497 4573 17509 4607
rect 17543 4573 17555 4607
rect 17497 4567 17555 4573
rect 14700 4508 15700 4536
rect 14700 4496 14706 4508
rect 17034 4496 17040 4548
rect 17092 4545 17098 4548
rect 17092 4536 17104 4545
rect 17092 4508 17137 4536
rect 17092 4499 17104 4508
rect 17092 4496 17098 4499
rect 10980 4440 12434 4468
rect 12710 4428 12716 4480
rect 12768 4428 12774 4480
rect 13446 4428 13452 4480
rect 13504 4468 13510 4480
rect 14366 4468 14372 4480
rect 13504 4440 14372 4468
rect 13504 4428 13510 4440
rect 14366 4428 14372 4440
rect 14424 4428 14430 4480
rect 15473 4471 15531 4477
rect 15473 4437 15485 4471
rect 15519 4468 15531 4471
rect 15562 4468 15568 4480
rect 15519 4440 15568 4468
rect 15519 4437 15531 4440
rect 15473 4431 15531 4437
rect 15562 4428 15568 4440
rect 15620 4428 15626 4480
rect 15654 4428 15660 4480
rect 15712 4468 15718 4480
rect 15933 4471 15991 4477
rect 15933 4468 15945 4471
rect 15712 4440 15945 4468
rect 15712 4428 15718 4440
rect 15933 4437 15945 4440
rect 15979 4437 15991 4471
rect 15933 4431 15991 4437
rect 1104 4378 18124 4400
rect 1104 4326 3737 4378
rect 3789 4326 3801 4378
rect 3853 4326 3865 4378
rect 3917 4326 3929 4378
rect 3981 4326 3993 4378
rect 4045 4326 7992 4378
rect 8044 4326 8056 4378
rect 8108 4326 8120 4378
rect 8172 4326 8184 4378
rect 8236 4326 8248 4378
rect 8300 4326 12247 4378
rect 12299 4326 12311 4378
rect 12363 4326 12375 4378
rect 12427 4326 12439 4378
rect 12491 4326 12503 4378
rect 12555 4326 16502 4378
rect 16554 4326 16566 4378
rect 16618 4326 16630 4378
rect 16682 4326 16694 4378
rect 16746 4326 16758 4378
rect 16810 4326 18124 4378
rect 1104 4304 18124 4326
rect 7374 4224 7380 4276
rect 7432 4264 7438 4276
rect 9858 4264 9864 4276
rect 7432 4236 9864 4264
rect 7432 4224 7438 4236
rect 9858 4224 9864 4236
rect 9916 4224 9922 4276
rect 11422 4224 11428 4276
rect 11480 4264 11486 4276
rect 11701 4267 11759 4273
rect 11701 4264 11713 4267
rect 11480 4236 11713 4264
rect 11480 4224 11486 4236
rect 11701 4233 11713 4236
rect 11747 4233 11759 4267
rect 11701 4227 11759 4233
rect 12069 4267 12127 4273
rect 12069 4233 12081 4267
rect 12115 4264 12127 4267
rect 12710 4264 12716 4276
rect 12115 4236 12716 4264
rect 12115 4233 12127 4236
rect 12069 4227 12127 4233
rect 12710 4224 12716 4236
rect 12768 4224 12774 4276
rect 13538 4224 13544 4276
rect 13596 4264 13602 4276
rect 13596 4236 14504 4264
rect 13596 4224 13602 4236
rect 6733 4199 6791 4205
rect 6733 4165 6745 4199
rect 6779 4196 6791 4199
rect 7193 4199 7251 4205
rect 7193 4196 7205 4199
rect 6779 4168 7205 4196
rect 6779 4165 6791 4168
rect 6733 4159 6791 4165
rect 7193 4165 7205 4168
rect 7239 4165 7251 4199
rect 14476 4196 14504 4236
rect 14550 4224 14556 4276
rect 14608 4264 14614 4276
rect 14645 4267 14703 4273
rect 14645 4264 14657 4267
rect 14608 4236 14657 4264
rect 14608 4224 14614 4236
rect 14645 4233 14657 4236
rect 14691 4233 14703 4267
rect 14645 4227 14703 4233
rect 15378 4224 15384 4276
rect 15436 4264 15442 4276
rect 15838 4264 15844 4276
rect 15436 4236 15844 4264
rect 15436 4224 15442 4236
rect 15838 4224 15844 4236
rect 15896 4224 15902 4276
rect 15470 4196 15476 4208
rect 14476 4168 15476 4196
rect 7193 4159 7251 4165
rect 15470 4156 15476 4168
rect 15528 4156 15534 4208
rect 15565 4199 15623 4205
rect 15565 4165 15577 4199
rect 15611 4196 15623 4199
rect 16390 4196 16396 4208
rect 15611 4168 16396 4196
rect 15611 4165 15623 4168
rect 15565 4159 15623 4165
rect 16390 4156 16396 4168
rect 16448 4156 16454 4208
rect 4982 4088 4988 4140
rect 5040 4128 5046 4140
rect 6825 4131 6883 4137
rect 6825 4128 6837 4131
rect 5040 4100 6837 4128
rect 5040 4088 5046 4100
rect 6825 4097 6837 4100
rect 6871 4097 6883 4131
rect 6825 4091 6883 4097
rect 7742 4088 7748 4140
rect 7800 4088 7806 4140
rect 9766 4088 9772 4140
rect 9824 4128 9830 4140
rect 9950 4128 9956 4140
rect 9824 4100 9956 4128
rect 9824 4088 9830 4100
rect 9950 4088 9956 4100
rect 10008 4128 10014 4140
rect 10505 4131 10563 4137
rect 10505 4128 10517 4131
rect 10008 4100 10517 4128
rect 10008 4088 10014 4100
rect 10505 4097 10517 4100
rect 10551 4097 10563 4131
rect 10505 4091 10563 4097
rect 10962 4088 10968 4140
rect 11020 4128 11026 4140
rect 11020 4100 12296 4128
rect 11020 4088 11026 4100
rect 5534 4020 5540 4072
rect 5592 4060 5598 4072
rect 5813 4063 5871 4069
rect 5813 4060 5825 4063
rect 5592 4032 5825 4060
rect 5592 4020 5598 4032
rect 5813 4029 5825 4032
rect 5859 4029 5871 4063
rect 5813 4023 5871 4029
rect 7009 4063 7067 4069
rect 7009 4029 7021 4063
rect 7055 4060 7067 4063
rect 8757 4063 8815 4069
rect 7055 4032 8524 4060
rect 7055 4029 7067 4032
rect 7009 4023 7067 4029
rect 5828 3992 5856 4023
rect 6730 3992 6736 4004
rect 5828 3964 6736 3992
rect 6730 3952 6736 3964
rect 6788 3992 6794 4004
rect 7190 3992 7196 4004
rect 6788 3964 7196 3992
rect 6788 3952 6794 3964
rect 7190 3952 7196 3964
rect 7248 3952 7254 4004
rect 4890 3884 4896 3936
rect 4948 3924 4954 3936
rect 5261 3927 5319 3933
rect 5261 3924 5273 3927
rect 4948 3896 5273 3924
rect 4948 3884 4954 3896
rect 5261 3893 5273 3896
rect 5307 3893 5319 3927
rect 5261 3887 5319 3893
rect 5810 3884 5816 3936
rect 5868 3924 5874 3936
rect 6365 3927 6423 3933
rect 6365 3924 6377 3927
rect 5868 3896 6377 3924
rect 5868 3884 5874 3896
rect 6365 3893 6377 3896
rect 6411 3893 6423 3927
rect 6365 3887 6423 3893
rect 8113 3927 8171 3933
rect 8113 3893 8125 3927
rect 8159 3924 8171 3927
rect 8386 3924 8392 3936
rect 8159 3896 8392 3924
rect 8159 3893 8171 3896
rect 8113 3887 8171 3893
rect 8386 3884 8392 3896
rect 8444 3884 8450 3936
rect 8496 3924 8524 4032
rect 8757 4029 8769 4063
rect 8803 4060 8815 4063
rect 9674 4060 9680 4072
rect 8803 4032 9680 4060
rect 8803 4029 8815 4032
rect 8757 4023 8815 4029
rect 9674 4020 9680 4032
rect 9732 4060 9738 4072
rect 10134 4060 10140 4072
rect 9732 4032 10140 4060
rect 9732 4020 9738 4032
rect 10134 4020 10140 4032
rect 10192 4020 10198 4072
rect 12268 4069 12296 4100
rect 12710 4088 12716 4140
rect 12768 4088 12774 4140
rect 12802 4088 12808 4140
rect 12860 4088 12866 4140
rect 13722 4088 13728 4140
rect 13780 4088 13786 4140
rect 13814 4088 13820 4140
rect 13872 4137 13878 4140
rect 13872 4131 13900 4137
rect 13888 4097 13900 4131
rect 13872 4091 13900 4097
rect 13872 4088 13878 4091
rect 13998 4088 14004 4140
rect 14056 4088 14062 4140
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 15746 4088 15752 4140
rect 15804 4128 15810 4140
rect 15841 4131 15899 4137
rect 15841 4128 15853 4131
rect 15804 4100 15853 4128
rect 15804 4088 15810 4100
rect 15841 4097 15853 4100
rect 15887 4097 15899 4131
rect 15841 4091 15899 4097
rect 16298 4088 16304 4140
rect 16356 4128 16362 4140
rect 16945 4131 17003 4137
rect 16945 4128 16957 4131
rect 16356 4100 16957 4128
rect 16356 4088 16362 4100
rect 16945 4097 16957 4100
rect 16991 4097 17003 4131
rect 16945 4091 17003 4097
rect 17494 4088 17500 4140
rect 17552 4088 17558 4140
rect 12161 4063 12219 4069
rect 12161 4029 12173 4063
rect 12207 4029 12219 4063
rect 12161 4023 12219 4029
rect 12253 4063 12311 4069
rect 12253 4029 12265 4063
rect 12299 4029 12311 4063
rect 12253 4023 12311 4029
rect 12989 4063 13047 4069
rect 12989 4029 13001 4063
rect 13035 4060 13047 4063
rect 13078 4060 13084 4072
rect 13035 4032 13084 4060
rect 13035 4029 13047 4032
rect 12989 4023 13047 4029
rect 8662 3952 8668 4004
rect 8720 3992 8726 4004
rect 11238 3992 11244 4004
rect 8720 3964 11244 3992
rect 8720 3952 8726 3964
rect 11238 3952 11244 3964
rect 11296 3952 11302 4004
rect 12176 3992 12204 4023
rect 13078 4020 13084 4032
rect 13136 4020 13142 4072
rect 13446 4020 13452 4072
rect 13504 4020 13510 4072
rect 15654 4020 15660 4072
rect 15712 4060 15718 4072
rect 16393 4063 16451 4069
rect 16393 4060 16405 4063
rect 15712 4032 16405 4060
rect 15712 4020 15718 4032
rect 16393 4029 16405 4032
rect 16439 4029 16451 4063
rect 16393 4023 16451 4029
rect 12434 3992 12440 4004
rect 12176 3964 12440 3992
rect 12434 3952 12440 3964
rect 12492 3992 12498 4004
rect 12492 3964 13584 3992
rect 12492 3952 12498 3964
rect 10134 3924 10140 3936
rect 8496 3896 10140 3924
rect 10134 3884 10140 3896
rect 10192 3924 10198 3936
rect 10686 3924 10692 3936
rect 10192 3896 10692 3924
rect 10192 3884 10198 3896
rect 10686 3884 10692 3896
rect 10744 3884 10750 3936
rect 10962 3884 10968 3936
rect 11020 3924 11026 3936
rect 11149 3927 11207 3933
rect 11149 3924 11161 3927
rect 11020 3896 11161 3924
rect 11020 3884 11026 3896
rect 11149 3893 11161 3896
rect 11195 3893 11207 3927
rect 11149 3887 11207 3893
rect 11974 3884 11980 3936
rect 12032 3924 12038 3936
rect 12529 3927 12587 3933
rect 12529 3924 12541 3927
rect 12032 3896 12541 3924
rect 12032 3884 12038 3896
rect 12529 3893 12541 3896
rect 12575 3893 12587 3927
rect 13556 3924 13584 3964
rect 15286 3924 15292 3936
rect 13556 3896 15292 3924
rect 12529 3887 12587 3893
rect 15286 3884 15292 3896
rect 15344 3884 15350 3936
rect 1104 3834 18124 3856
rect 1104 3782 3077 3834
rect 3129 3782 3141 3834
rect 3193 3782 3205 3834
rect 3257 3782 3269 3834
rect 3321 3782 3333 3834
rect 3385 3782 7332 3834
rect 7384 3782 7396 3834
rect 7448 3782 7460 3834
rect 7512 3782 7524 3834
rect 7576 3782 7588 3834
rect 7640 3782 11587 3834
rect 11639 3782 11651 3834
rect 11703 3782 11715 3834
rect 11767 3782 11779 3834
rect 11831 3782 11843 3834
rect 11895 3782 15842 3834
rect 15894 3782 15906 3834
rect 15958 3782 15970 3834
rect 16022 3782 16034 3834
rect 16086 3782 16098 3834
rect 16150 3782 18124 3834
rect 1104 3760 18124 3782
rect 6733 3723 6791 3729
rect 6733 3689 6745 3723
rect 6779 3720 6791 3723
rect 7006 3720 7012 3732
rect 6779 3692 7012 3720
rect 6779 3689 6791 3692
rect 6733 3683 6791 3689
rect 7006 3680 7012 3692
rect 7064 3680 7070 3732
rect 7098 3680 7104 3732
rect 7156 3720 7162 3732
rect 7156 3692 15424 3720
rect 7156 3680 7162 3692
rect 4525 3655 4583 3661
rect 4525 3621 4537 3655
rect 4571 3621 4583 3655
rect 4525 3615 4583 3621
rect 8757 3655 8815 3661
rect 8757 3621 8769 3655
rect 8803 3621 8815 3655
rect 8757 3615 8815 3621
rect 4433 3519 4491 3525
rect 4433 3485 4445 3519
rect 4479 3516 4491 3519
rect 4540 3516 4568 3615
rect 4982 3544 4988 3596
rect 5040 3544 5046 3596
rect 5169 3587 5227 3593
rect 5169 3553 5181 3587
rect 5215 3584 5227 3587
rect 5215 3556 5488 3584
rect 5215 3553 5227 3556
rect 5169 3547 5227 3553
rect 4479 3488 4568 3516
rect 4479 3485 4491 3488
rect 4433 3479 4491 3485
rect 4890 3476 4896 3528
rect 4948 3476 4954 3528
rect 5353 3519 5411 3525
rect 5353 3485 5365 3519
rect 5399 3485 5411 3519
rect 5460 3516 5488 3556
rect 7098 3544 7104 3596
rect 7156 3544 7162 3596
rect 8205 3587 8263 3593
rect 8205 3553 8217 3587
rect 8251 3584 8263 3587
rect 8662 3584 8668 3596
rect 8251 3556 8668 3584
rect 8251 3553 8263 3556
rect 8205 3547 8263 3553
rect 5460 3488 5764 3516
rect 5353 3479 5411 3485
rect 4154 3408 4160 3460
rect 4212 3448 4218 3460
rect 5368 3448 5396 3479
rect 5626 3457 5632 3460
rect 4212 3420 5396 3448
rect 4212 3408 4218 3420
rect 5620 3411 5632 3457
rect 5626 3408 5632 3411
rect 5684 3408 5690 3460
rect 5736 3448 5764 3488
rect 7190 3476 7196 3528
rect 7248 3516 7254 3528
rect 7285 3519 7343 3525
rect 7285 3516 7297 3519
rect 7248 3488 7297 3516
rect 7248 3476 7254 3488
rect 7285 3485 7297 3488
rect 7331 3485 7343 3519
rect 7285 3479 7343 3485
rect 8220 3448 8248 3547
rect 8662 3544 8668 3556
rect 8720 3544 8726 3596
rect 8386 3476 8392 3528
rect 8444 3476 8450 3528
rect 8772 3516 8800 3615
rect 10594 3612 10600 3664
rect 10652 3612 10658 3664
rect 11072 3652 11100 3692
rect 11072 3624 11192 3652
rect 9324 3556 9812 3584
rect 9125 3519 9183 3525
rect 9125 3516 9137 3519
rect 8772 3488 9137 3516
rect 9125 3485 9137 3488
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 5736 3420 8248 3448
rect 8297 3451 8355 3457
rect 8297 3417 8309 3451
rect 8343 3448 8355 3451
rect 8846 3448 8852 3460
rect 8343 3420 8852 3448
rect 8343 3417 8355 3420
rect 8297 3411 8355 3417
rect 8846 3408 8852 3420
rect 8904 3448 8910 3460
rect 9324 3448 9352 3556
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3516 9459 3519
rect 9447 3488 9536 3516
rect 9447 3485 9459 3488
rect 9401 3479 9459 3485
rect 8904 3420 9352 3448
rect 8904 3408 8910 3420
rect 4246 3340 4252 3392
rect 4304 3340 4310 3392
rect 4982 3340 4988 3392
rect 5040 3380 5046 3392
rect 7193 3383 7251 3389
rect 7193 3380 7205 3383
rect 5040 3352 7205 3380
rect 5040 3340 5046 3352
rect 7193 3349 7205 3352
rect 7239 3349 7251 3383
rect 7193 3343 7251 3349
rect 7653 3383 7711 3389
rect 7653 3349 7665 3383
rect 7699 3380 7711 3383
rect 7742 3380 7748 3392
rect 7699 3352 7748 3380
rect 7699 3349 7711 3352
rect 7653 3343 7711 3349
rect 7742 3340 7748 3352
rect 7800 3340 7806 3392
rect 8938 3340 8944 3392
rect 8996 3340 9002 3392
rect 9217 3383 9275 3389
rect 9217 3349 9229 3383
rect 9263 3380 9275 3383
rect 9306 3380 9312 3392
rect 9263 3352 9312 3380
rect 9263 3349 9275 3352
rect 9217 3343 9275 3349
rect 9306 3340 9312 3352
rect 9364 3340 9370 3392
rect 9508 3389 9536 3488
rect 9493 3383 9551 3389
rect 9493 3349 9505 3383
rect 9539 3349 9551 3383
rect 9784 3380 9812 3556
rect 10134 3544 10140 3596
rect 10192 3544 10198 3596
rect 10410 3544 10416 3596
rect 10468 3584 10474 3596
rect 11164 3593 11192 3624
rect 12710 3612 12716 3664
rect 12768 3652 12774 3664
rect 12989 3655 13047 3661
rect 12989 3652 13001 3655
rect 12768 3624 13001 3652
rect 12768 3612 12774 3624
rect 12989 3621 13001 3624
rect 13035 3621 13047 3655
rect 12989 3615 13047 3621
rect 14829 3655 14887 3661
rect 14829 3621 14841 3655
rect 14875 3621 14887 3655
rect 14829 3615 14887 3621
rect 11149 3587 11207 3593
rect 10468 3556 11100 3584
rect 10468 3544 10474 3556
rect 10962 3476 10968 3528
rect 11020 3476 11026 3528
rect 11072 3516 11100 3556
rect 11149 3553 11161 3587
rect 11195 3553 11207 3587
rect 11149 3547 11207 3553
rect 11238 3544 11244 3596
rect 11296 3584 11302 3596
rect 12345 3587 12403 3593
rect 12345 3584 12357 3587
rect 11296 3556 12357 3584
rect 11296 3544 11302 3556
rect 12345 3553 12357 3556
rect 12391 3553 12403 3587
rect 12345 3547 12403 3553
rect 12434 3544 12440 3596
rect 12492 3584 12498 3596
rect 12529 3587 12587 3593
rect 12529 3584 12541 3587
rect 12492 3556 12541 3584
rect 12492 3544 12498 3556
rect 12529 3553 12541 3556
rect 12575 3553 12587 3587
rect 12529 3547 12587 3553
rect 13722 3544 13728 3596
rect 13780 3544 13786 3596
rect 11977 3519 12035 3525
rect 11977 3516 11989 3519
rect 11072 3488 11989 3516
rect 11977 3485 11989 3488
rect 12023 3485 12035 3519
rect 13538 3516 13544 3528
rect 11977 3479 12035 3485
rect 12406 3488 13544 3516
rect 9861 3451 9919 3457
rect 9861 3417 9873 3451
rect 9907 3448 9919 3451
rect 11425 3451 11483 3457
rect 11425 3448 11437 3451
rect 9907 3420 11437 3448
rect 9907 3417 9919 3420
rect 9861 3411 9919 3417
rect 11425 3417 11437 3420
rect 11471 3417 11483 3451
rect 11425 3411 11483 3417
rect 9953 3383 10011 3389
rect 9953 3380 9965 3383
rect 9784 3352 9965 3380
rect 9493 3343 9551 3349
rect 9953 3349 9965 3352
rect 9999 3380 10011 3383
rect 11057 3383 11115 3389
rect 11057 3380 11069 3383
rect 9999 3352 11069 3380
rect 9999 3349 10011 3352
rect 9953 3343 10011 3349
rect 11057 3349 11069 3352
rect 11103 3380 11115 3383
rect 12406 3380 12434 3488
rect 13538 3476 13544 3488
rect 13596 3476 13602 3528
rect 14090 3476 14096 3528
rect 14148 3476 14154 3528
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3516 14611 3519
rect 14844 3516 14872 3615
rect 15286 3544 15292 3596
rect 15344 3544 15350 3596
rect 15396 3593 15424 3692
rect 15381 3587 15439 3593
rect 15381 3553 15393 3587
rect 15427 3553 15439 3587
rect 15381 3547 15439 3553
rect 16022 3516 16028 3528
rect 14599 3488 14872 3516
rect 14936 3488 16028 3516
rect 14599 3485 14611 3488
rect 14553 3479 14611 3485
rect 12621 3451 12679 3457
rect 12621 3417 12633 3451
rect 12667 3448 12679 3451
rect 13081 3451 13139 3457
rect 13081 3448 13093 3451
rect 12667 3420 13093 3448
rect 12667 3417 12679 3420
rect 12621 3411 12679 3417
rect 13081 3417 13093 3420
rect 13127 3417 13139 3451
rect 13081 3411 13139 3417
rect 13170 3408 13176 3460
rect 13228 3448 13234 3460
rect 14936 3448 14964 3488
rect 16022 3476 16028 3488
rect 16080 3516 16086 3528
rect 16209 3519 16267 3525
rect 16209 3516 16221 3519
rect 16080 3488 16221 3516
rect 16080 3476 16086 3488
rect 16209 3485 16221 3488
rect 16255 3485 16267 3519
rect 16209 3479 16267 3485
rect 13228 3420 14964 3448
rect 15197 3451 15255 3457
rect 13228 3408 13234 3420
rect 15197 3417 15209 3451
rect 15243 3448 15255 3451
rect 15657 3451 15715 3457
rect 15657 3448 15669 3451
rect 15243 3420 15669 3448
rect 15243 3417 15255 3420
rect 15197 3411 15255 3417
rect 15657 3417 15669 3420
rect 15703 3417 15715 3451
rect 15657 3411 15715 3417
rect 17678 3408 17684 3460
rect 17736 3408 17742 3460
rect 11103 3352 12434 3380
rect 11103 3349 11115 3352
rect 11057 3343 11115 3349
rect 14274 3340 14280 3392
rect 14332 3340 14338 3392
rect 14734 3340 14740 3392
rect 14792 3340 14798 3392
rect 14918 3340 14924 3392
rect 14976 3380 14982 3392
rect 15286 3380 15292 3392
rect 14976 3352 15292 3380
rect 14976 3340 14982 3352
rect 15286 3340 15292 3352
rect 15344 3380 15350 3392
rect 17589 3383 17647 3389
rect 17589 3380 17601 3383
rect 15344 3352 17601 3380
rect 15344 3340 15350 3352
rect 17589 3349 17601 3352
rect 17635 3349 17647 3383
rect 17589 3343 17647 3349
rect 1104 3290 18124 3312
rect 1104 3238 3737 3290
rect 3789 3238 3801 3290
rect 3853 3238 3865 3290
rect 3917 3238 3929 3290
rect 3981 3238 3993 3290
rect 4045 3238 7992 3290
rect 8044 3238 8056 3290
rect 8108 3238 8120 3290
rect 8172 3238 8184 3290
rect 8236 3238 8248 3290
rect 8300 3238 12247 3290
rect 12299 3238 12311 3290
rect 12363 3238 12375 3290
rect 12427 3238 12439 3290
rect 12491 3238 12503 3290
rect 12555 3238 16502 3290
rect 16554 3238 16566 3290
rect 16618 3238 16630 3290
rect 16682 3238 16694 3290
rect 16746 3238 16758 3290
rect 16810 3238 18124 3290
rect 1104 3216 18124 3238
rect 5534 3136 5540 3188
rect 5592 3136 5598 3188
rect 5626 3136 5632 3188
rect 5684 3136 5690 3188
rect 6365 3179 6423 3185
rect 6365 3145 6377 3179
rect 6411 3176 6423 3179
rect 6822 3176 6828 3188
rect 6411 3148 6828 3176
rect 6411 3145 6423 3148
rect 6365 3139 6423 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 9217 3179 9275 3185
rect 9217 3145 9229 3179
rect 9263 3176 9275 3179
rect 9674 3176 9680 3188
rect 9263 3148 9680 3176
rect 9263 3145 9275 3148
rect 9217 3139 9275 3145
rect 9674 3136 9680 3148
rect 9732 3136 9738 3188
rect 9861 3179 9919 3185
rect 9861 3145 9873 3179
rect 9907 3145 9919 3179
rect 9861 3139 9919 3145
rect 4246 3068 4252 3120
rect 4304 3108 4310 3120
rect 4402 3111 4460 3117
rect 4402 3108 4414 3111
rect 4304 3080 4414 3108
rect 4304 3068 4310 3080
rect 4402 3077 4414 3080
rect 4448 3077 4460 3111
rect 4402 3071 4460 3077
rect 8104 3111 8162 3117
rect 8104 3077 8116 3111
rect 8150 3108 8162 3111
rect 8938 3108 8944 3120
rect 8150 3080 8944 3108
rect 8150 3077 8162 3080
rect 8104 3071 8162 3077
rect 8938 3068 8944 3080
rect 8996 3068 9002 3120
rect 9876 3108 9904 3139
rect 9950 3136 9956 3188
rect 10008 3136 10014 3188
rect 12802 3136 12808 3188
rect 12860 3176 12866 3188
rect 13170 3176 13176 3188
rect 12860 3148 13176 3176
rect 12860 3136 12866 3148
rect 13170 3136 13176 3148
rect 13228 3136 13234 3188
rect 16022 3136 16028 3188
rect 16080 3136 16086 3188
rect 11066 3111 11124 3117
rect 11066 3108 11078 3111
rect 9876 3080 11078 3108
rect 11066 3077 11078 3080
rect 11112 3077 11124 3111
rect 12618 3108 12624 3120
rect 11066 3071 11124 3077
rect 11716 3080 12624 3108
rect 4154 3000 4160 3052
rect 4212 3000 4218 3052
rect 5810 3000 5816 3052
rect 5868 3000 5874 3052
rect 7489 3043 7547 3049
rect 7489 3009 7501 3043
rect 7535 3040 7547 3043
rect 7650 3040 7656 3052
rect 7535 3012 7656 3040
rect 7535 3009 7547 3012
rect 7489 3003 7547 3009
rect 7650 3000 7656 3012
rect 7708 3000 7714 3052
rect 7745 3043 7803 3049
rect 7745 3009 7757 3043
rect 7791 3040 7803 3043
rect 7837 3043 7895 3049
rect 7837 3040 7849 3043
rect 7791 3012 7849 3040
rect 7791 3009 7803 3012
rect 7745 3003 7803 3009
rect 7837 3009 7849 3012
rect 7883 3040 7895 3043
rect 7926 3040 7932 3052
rect 7883 3012 7932 3040
rect 7883 3009 7895 3012
rect 7837 3003 7895 3009
rect 7926 3000 7932 3012
rect 7984 3000 7990 3052
rect 9030 3000 9036 3052
rect 9088 3040 9094 3052
rect 9401 3043 9459 3049
rect 9401 3040 9413 3043
rect 9088 3012 9413 3040
rect 9088 3000 9094 3012
rect 9401 3009 9413 3012
rect 9447 3009 9459 3043
rect 9401 3003 9459 3009
rect 9677 3043 9735 3049
rect 9677 3009 9689 3043
rect 9723 3040 9735 3043
rect 10594 3040 10600 3052
rect 9723 3012 10600 3040
rect 9723 3009 9735 3012
rect 9677 3003 9735 3009
rect 10594 3000 10600 3012
rect 10652 3000 10658 3052
rect 11716 3049 11744 3080
rect 12618 3068 12624 3080
rect 12676 3108 12682 3120
rect 12676 3080 14596 3108
rect 12676 3068 12682 3080
rect 11974 3049 11980 3052
rect 11333 3043 11391 3049
rect 11333 3009 11345 3043
rect 11379 3040 11391 3043
rect 11701 3043 11759 3049
rect 11701 3040 11713 3043
rect 11379 3012 11713 3040
rect 11379 3009 11391 3012
rect 11333 3003 11391 3009
rect 11701 3009 11713 3012
rect 11747 3009 11759 3043
rect 11968 3040 11980 3049
rect 11935 3012 11980 3040
rect 11701 3003 11759 3009
rect 11968 3003 11980 3012
rect 11974 3000 11980 3003
rect 12032 3000 12038 3052
rect 14274 3000 14280 3052
rect 14332 3049 14338 3052
rect 14568 3049 14596 3080
rect 14734 3068 14740 3120
rect 14792 3108 14798 3120
rect 14890 3111 14948 3117
rect 14890 3108 14902 3111
rect 14792 3080 14902 3108
rect 14792 3068 14798 3080
rect 14890 3077 14902 3080
rect 14936 3077 14948 3111
rect 14890 3071 14948 3077
rect 14332 3040 14344 3049
rect 14553 3043 14611 3049
rect 14332 3012 14377 3040
rect 14332 3003 14344 3012
rect 14553 3009 14565 3043
rect 14599 3009 14611 3043
rect 14553 3003 14611 3009
rect 14332 3000 14338 3003
rect 14642 3000 14648 3052
rect 14700 3000 14706 3052
rect 9398 2796 9404 2848
rect 9456 2836 9462 2848
rect 9493 2839 9551 2845
rect 9493 2836 9505 2839
rect 9456 2808 9505 2836
rect 9456 2796 9462 2808
rect 9493 2805 9505 2808
rect 9539 2805 9551 2839
rect 9493 2799 9551 2805
rect 13081 2839 13139 2845
rect 13081 2805 13093 2839
rect 13127 2836 13139 2839
rect 13630 2836 13636 2848
rect 13127 2808 13636 2836
rect 13127 2805 13139 2808
rect 13081 2799 13139 2805
rect 13630 2796 13636 2808
rect 13688 2796 13694 2848
rect 1104 2746 18124 2768
rect 1104 2694 3077 2746
rect 3129 2694 3141 2746
rect 3193 2694 3205 2746
rect 3257 2694 3269 2746
rect 3321 2694 3333 2746
rect 3385 2694 7332 2746
rect 7384 2694 7396 2746
rect 7448 2694 7460 2746
rect 7512 2694 7524 2746
rect 7576 2694 7588 2746
rect 7640 2694 11587 2746
rect 11639 2694 11651 2746
rect 11703 2694 11715 2746
rect 11767 2694 11779 2746
rect 11831 2694 11843 2746
rect 11895 2694 15842 2746
rect 15894 2694 15906 2746
rect 15958 2694 15970 2746
rect 16022 2694 16034 2746
rect 16086 2694 16098 2746
rect 16150 2694 18124 2746
rect 1104 2672 18124 2694
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7561 2635 7619 2641
rect 7561 2632 7573 2635
rect 7248 2604 7573 2632
rect 7248 2592 7254 2604
rect 7561 2601 7573 2604
rect 7607 2601 7619 2635
rect 7561 2595 7619 2601
rect 7650 2592 7656 2644
rect 7708 2592 7714 2644
rect 10410 2592 10416 2644
rect 10468 2592 10474 2644
rect 14090 2592 14096 2644
rect 14148 2592 14154 2644
rect 4249 2567 4307 2573
rect 4249 2533 4261 2567
rect 4295 2564 4307 2567
rect 4982 2564 4988 2576
rect 4295 2536 4988 2564
rect 4295 2533 4307 2536
rect 4249 2527 4307 2533
rect 4982 2524 4988 2536
rect 5040 2524 5046 2576
rect 11606 2524 11612 2576
rect 11664 2564 11670 2576
rect 12989 2567 13047 2573
rect 12989 2564 13001 2567
rect 11664 2536 13001 2564
rect 11664 2524 11670 2536
rect 12989 2533 13001 2536
rect 13035 2533 13047 2567
rect 12989 2527 13047 2533
rect 13449 2567 13507 2573
rect 13449 2533 13461 2567
rect 13495 2564 13507 2567
rect 13538 2564 13544 2576
rect 13495 2536 13544 2564
rect 13495 2533 13507 2536
rect 13449 2527 13507 2533
rect 13538 2524 13544 2536
rect 13596 2524 13602 2576
rect 14918 2564 14924 2576
rect 14568 2536 14924 2564
rect 6822 2456 6828 2508
rect 6880 2496 6886 2508
rect 6917 2499 6975 2505
rect 6917 2496 6929 2499
rect 6880 2468 6929 2496
rect 6880 2456 6886 2468
rect 6917 2465 6929 2468
rect 6963 2465 6975 2499
rect 6917 2459 6975 2465
rect 7926 2456 7932 2508
rect 7984 2496 7990 2508
rect 9033 2499 9091 2505
rect 9033 2496 9045 2499
rect 7984 2468 9045 2496
rect 7984 2456 7990 2468
rect 9033 2465 9045 2468
rect 9079 2465 9091 2499
rect 9033 2459 9091 2465
rect 10781 2499 10839 2505
rect 10781 2465 10793 2499
rect 10827 2496 10839 2499
rect 10870 2496 10876 2508
rect 10827 2468 10876 2496
rect 10827 2465 10839 2468
rect 10781 2459 10839 2465
rect 10870 2456 10876 2468
rect 10928 2456 10934 2508
rect 11793 2499 11851 2505
rect 11793 2465 11805 2499
rect 11839 2496 11851 2499
rect 12066 2496 12072 2508
rect 11839 2468 12072 2496
rect 11839 2465 11851 2468
rect 11793 2459 11851 2465
rect 12066 2456 12072 2468
rect 12124 2456 12130 2508
rect 14568 2505 14596 2536
rect 14918 2524 14924 2536
rect 14976 2524 14982 2576
rect 14553 2499 14611 2505
rect 14553 2465 14565 2499
rect 14599 2465 14611 2499
rect 14553 2459 14611 2465
rect 14642 2456 14648 2508
rect 14700 2456 14706 2508
rect 5905 2431 5963 2437
rect 5905 2397 5917 2431
rect 5951 2428 5963 2431
rect 6086 2428 6092 2440
rect 5951 2400 6092 2428
rect 5951 2397 5963 2400
rect 5905 2391 5963 2397
rect 6086 2388 6092 2400
rect 6144 2388 6150 2440
rect 6270 2388 6276 2440
rect 6328 2428 6334 2440
rect 6549 2431 6607 2437
rect 6549 2428 6561 2431
rect 6328 2400 6561 2428
rect 6328 2388 6334 2400
rect 6549 2397 6561 2400
rect 6595 2397 6607 2431
rect 6549 2391 6607 2397
rect 7834 2388 7840 2440
rect 7892 2388 7898 2440
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 9306 2437 9312 2440
rect 8757 2431 8815 2437
rect 8757 2397 8769 2431
rect 8803 2397 8815 2431
rect 9300 2428 9312 2437
rect 9267 2400 9312 2428
rect 8757 2391 8815 2397
rect 9300 2391 9312 2400
rect 4062 2320 4068 2372
rect 4120 2320 4126 2372
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 8772 2360 8800 2391
rect 9306 2388 9312 2391
rect 9364 2388 9370 2440
rect 10318 2388 10324 2440
rect 10376 2428 10382 2440
rect 10505 2431 10563 2437
rect 10505 2428 10517 2431
rect 10376 2400 10517 2428
rect 10376 2388 10382 2400
rect 10505 2397 10517 2400
rect 10551 2397 10563 2431
rect 10505 2391 10563 2397
rect 11517 2431 11575 2437
rect 11517 2397 11529 2431
rect 11563 2397 11575 2431
rect 11517 2391 11575 2397
rect 12437 2431 12495 2437
rect 12437 2397 12449 2431
rect 12483 2428 12495 2431
rect 12710 2428 12716 2440
rect 12483 2400 12716 2428
rect 12483 2397 12495 2400
rect 12437 2391 12495 2397
rect 8444 2332 8800 2360
rect 8444 2320 8450 2332
rect 9674 2320 9680 2372
rect 9732 2360 9738 2372
rect 11532 2360 11560 2391
rect 12710 2388 12716 2400
rect 12768 2388 12774 2440
rect 12805 2431 12863 2437
rect 12805 2397 12817 2431
rect 12851 2428 12863 2431
rect 12894 2428 12900 2440
rect 12851 2400 12900 2428
rect 12851 2397 12863 2400
rect 12805 2391 12863 2397
rect 12894 2388 12900 2400
rect 12952 2388 12958 2440
rect 13170 2388 13176 2440
rect 13228 2428 13234 2440
rect 15473 2431 15531 2437
rect 15473 2428 15485 2431
rect 13228 2400 15485 2428
rect 13228 2388 13234 2400
rect 15473 2397 15485 2400
rect 15519 2397 15531 2431
rect 15473 2391 15531 2397
rect 9732 2332 11560 2360
rect 9732 2320 9738 2332
rect 12158 2320 12164 2372
rect 12216 2360 12222 2372
rect 13265 2363 13323 2369
rect 13265 2360 13277 2363
rect 12216 2332 13277 2360
rect 12216 2320 12222 2332
rect 13265 2329 13277 2332
rect 13311 2329 13323 2363
rect 13265 2323 13323 2329
rect 14461 2363 14519 2369
rect 14461 2329 14473 2363
rect 14507 2360 14519 2363
rect 14921 2363 14979 2369
rect 14921 2360 14933 2363
rect 14507 2332 14933 2360
rect 14507 2329 14519 2332
rect 14461 2323 14519 2329
rect 14921 2329 14933 2332
rect 14967 2329 14979 2363
rect 14921 2323 14979 2329
rect 6089 2295 6147 2301
rect 6089 2261 6101 2295
rect 6135 2292 6147 2295
rect 6454 2292 6460 2304
rect 6135 2264 6460 2292
rect 6135 2261 6147 2264
rect 6089 2255 6147 2261
rect 6454 2252 6460 2264
rect 6512 2252 6518 2304
rect 6733 2295 6791 2301
rect 6733 2261 6745 2295
rect 6779 2292 6791 2295
rect 7098 2292 7104 2304
rect 6779 2264 7104 2292
rect 6779 2261 6791 2264
rect 6733 2255 6791 2261
rect 7098 2252 7104 2264
rect 7156 2252 7162 2304
rect 10962 2252 10968 2304
rect 11020 2292 11026 2304
rect 12621 2295 12679 2301
rect 12621 2292 12633 2295
rect 11020 2264 12633 2292
rect 11020 2252 11026 2264
rect 12621 2261 12633 2264
rect 12667 2261 12679 2295
rect 12621 2255 12679 2261
rect 1104 2202 18124 2224
rect 1104 2150 3737 2202
rect 3789 2150 3801 2202
rect 3853 2150 3865 2202
rect 3917 2150 3929 2202
rect 3981 2150 3993 2202
rect 4045 2150 7992 2202
rect 8044 2150 8056 2202
rect 8108 2150 8120 2202
rect 8172 2150 8184 2202
rect 8236 2150 8248 2202
rect 8300 2150 12247 2202
rect 12299 2150 12311 2202
rect 12363 2150 12375 2202
rect 12427 2150 12439 2202
rect 12491 2150 12503 2202
rect 12555 2150 16502 2202
rect 16554 2150 16566 2202
rect 16618 2150 16630 2202
rect 16682 2150 16694 2202
rect 16746 2150 16758 2202
rect 16810 2150 18124 2202
rect 1104 2128 18124 2150
<< via1 >>
rect 3077 19014 3129 19066
rect 3141 19014 3193 19066
rect 3205 19014 3257 19066
rect 3269 19014 3321 19066
rect 3333 19014 3385 19066
rect 7332 19014 7384 19066
rect 7396 19014 7448 19066
rect 7460 19014 7512 19066
rect 7524 19014 7576 19066
rect 7588 19014 7640 19066
rect 11587 19014 11639 19066
rect 11651 19014 11703 19066
rect 11715 19014 11767 19066
rect 11779 19014 11831 19066
rect 11843 19014 11895 19066
rect 15842 19014 15894 19066
rect 15906 19014 15958 19066
rect 15970 19014 16022 19066
rect 16034 19014 16086 19066
rect 16098 19014 16150 19066
rect 10324 18912 10376 18964
rect 12624 18955 12676 18964
rect 12624 18921 12633 18955
rect 12633 18921 12667 18955
rect 12667 18921 12676 18955
rect 12624 18912 12676 18921
rect 7104 18751 7156 18760
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 7840 18708 7892 18760
rect 8576 18708 8628 18760
rect 9036 18708 9088 18760
rect 9312 18708 9364 18760
rect 10600 18708 10652 18760
rect 11152 18751 11204 18760
rect 11152 18717 11161 18751
rect 11161 18717 11195 18751
rect 11195 18717 11204 18751
rect 11152 18708 11204 18717
rect 12624 18708 12676 18760
rect 13084 18708 13136 18760
rect 13820 18751 13872 18760
rect 13820 18717 13829 18751
rect 13829 18717 13863 18751
rect 13863 18717 13872 18751
rect 13820 18708 13872 18717
rect 8484 18683 8536 18692
rect 8484 18649 8493 18683
rect 8493 18649 8527 18683
rect 8527 18649 8536 18683
rect 8484 18640 8536 18649
rect 9772 18683 9824 18692
rect 9772 18649 9781 18683
rect 9781 18649 9815 18683
rect 9815 18649 9824 18683
rect 9772 18640 9824 18649
rect 14096 18640 14148 18692
rect 6736 18572 6788 18624
rect 7656 18615 7708 18624
rect 7656 18581 7665 18615
rect 7665 18581 7699 18615
rect 7699 18581 7708 18615
rect 7656 18572 7708 18581
rect 7748 18615 7800 18624
rect 7748 18581 7757 18615
rect 7757 18581 7791 18615
rect 7791 18581 7800 18615
rect 7748 18572 7800 18581
rect 8944 18615 8996 18624
rect 8944 18581 8953 18615
rect 8953 18581 8987 18615
rect 8987 18581 8996 18615
rect 8944 18572 8996 18581
rect 9864 18572 9916 18624
rect 11336 18615 11388 18624
rect 11336 18581 11345 18615
rect 11345 18581 11379 18615
rect 11379 18581 11388 18615
rect 11336 18572 11388 18581
rect 11428 18572 11480 18624
rect 12900 18615 12952 18624
rect 12900 18581 12909 18615
rect 12909 18581 12943 18615
rect 12943 18581 12952 18615
rect 12900 18572 12952 18581
rect 13636 18615 13688 18624
rect 13636 18581 13645 18615
rect 13645 18581 13679 18615
rect 13679 18581 13688 18615
rect 13636 18572 13688 18581
rect 3737 18470 3789 18522
rect 3801 18470 3853 18522
rect 3865 18470 3917 18522
rect 3929 18470 3981 18522
rect 3993 18470 4045 18522
rect 7992 18470 8044 18522
rect 8056 18470 8108 18522
rect 8120 18470 8172 18522
rect 8184 18470 8236 18522
rect 8248 18470 8300 18522
rect 12247 18470 12299 18522
rect 12311 18470 12363 18522
rect 12375 18470 12427 18522
rect 12439 18470 12491 18522
rect 12503 18470 12555 18522
rect 16502 18470 16554 18522
rect 16566 18470 16618 18522
rect 16630 18470 16682 18522
rect 16694 18470 16746 18522
rect 16758 18470 16810 18522
rect 7656 18368 7708 18420
rect 9312 18411 9364 18420
rect 9312 18377 9321 18411
rect 9321 18377 9355 18411
rect 9355 18377 9364 18411
rect 9312 18368 9364 18377
rect 9680 18368 9732 18420
rect 10508 18368 10560 18420
rect 11980 18368 12032 18420
rect 13084 18411 13136 18420
rect 13084 18377 13093 18411
rect 13093 18377 13127 18411
rect 13127 18377 13136 18411
rect 13084 18368 13136 18377
rect 6736 18275 6788 18284
rect 6736 18241 6770 18275
rect 6770 18241 6788 18275
rect 6736 18232 6788 18241
rect 11060 18300 11112 18352
rect 10692 18232 10744 18284
rect 7748 18164 7800 18216
rect 11336 18164 11388 18216
rect 13636 18300 13688 18352
rect 15660 18275 15712 18284
rect 15660 18241 15669 18275
rect 15669 18241 15703 18275
rect 15703 18241 15712 18275
rect 15660 18232 15712 18241
rect 15016 18096 15068 18148
rect 8576 18028 8628 18080
rect 9496 18028 9548 18080
rect 12624 18028 12676 18080
rect 14740 18071 14792 18080
rect 14740 18037 14749 18071
rect 14749 18037 14783 18071
rect 14783 18037 14792 18071
rect 14740 18028 14792 18037
rect 15384 18028 15436 18080
rect 3077 17926 3129 17978
rect 3141 17926 3193 17978
rect 3205 17926 3257 17978
rect 3269 17926 3321 17978
rect 3333 17926 3385 17978
rect 7332 17926 7384 17978
rect 7396 17926 7448 17978
rect 7460 17926 7512 17978
rect 7524 17926 7576 17978
rect 7588 17926 7640 17978
rect 11587 17926 11639 17978
rect 11651 17926 11703 17978
rect 11715 17926 11767 17978
rect 11779 17926 11831 17978
rect 11843 17926 11895 17978
rect 15842 17926 15894 17978
rect 15906 17926 15958 17978
rect 15970 17926 16022 17978
rect 16034 17926 16086 17978
rect 16098 17926 16150 17978
rect 7104 17824 7156 17876
rect 7840 17824 7892 17876
rect 5172 17688 5224 17740
rect 8392 17756 8444 17808
rect 10140 17824 10192 17876
rect 10600 17824 10652 17876
rect 10692 17867 10744 17876
rect 10692 17833 10701 17867
rect 10701 17833 10735 17867
rect 10735 17833 10744 17867
rect 10692 17824 10744 17833
rect 11152 17824 11204 17876
rect 13820 17824 13872 17876
rect 4712 17663 4764 17672
rect 4712 17629 4721 17663
rect 4721 17629 4755 17663
rect 4755 17629 4764 17663
rect 4712 17620 4764 17629
rect 5080 17663 5132 17672
rect 5080 17629 5089 17663
rect 5089 17629 5123 17663
rect 5123 17629 5132 17663
rect 5080 17620 5132 17629
rect 5632 17663 5684 17672
rect 5632 17629 5641 17663
rect 5641 17629 5675 17663
rect 5675 17629 5684 17663
rect 5632 17620 5684 17629
rect 8576 17688 8628 17740
rect 8668 17731 8720 17740
rect 8668 17697 8677 17731
rect 8677 17697 8711 17731
rect 8711 17697 8720 17731
rect 8668 17688 8720 17697
rect 11520 17731 11572 17740
rect 4436 17552 4488 17604
rect 7656 17620 7708 17672
rect 7748 17620 7800 17672
rect 8944 17552 8996 17604
rect 10232 17552 10284 17604
rect 4160 17527 4212 17536
rect 4160 17493 4169 17527
rect 4169 17493 4203 17527
rect 4203 17493 4212 17527
rect 4160 17484 4212 17493
rect 4896 17527 4948 17536
rect 4896 17493 4905 17527
rect 4905 17493 4939 17527
rect 4939 17493 4948 17527
rect 4896 17484 4948 17493
rect 6000 17484 6052 17536
rect 8484 17527 8536 17536
rect 8484 17493 8493 17527
rect 8493 17493 8527 17527
rect 8527 17493 8536 17527
rect 8484 17484 8536 17493
rect 8576 17484 8628 17536
rect 11520 17697 11529 17731
rect 11529 17697 11563 17731
rect 11563 17697 11572 17731
rect 11520 17688 11572 17697
rect 12440 17756 12492 17808
rect 13176 17688 13228 17740
rect 16212 17688 16264 17740
rect 11428 17620 11480 17672
rect 12440 17620 12492 17672
rect 12900 17620 12952 17672
rect 14924 17620 14976 17672
rect 15384 17663 15436 17672
rect 15384 17629 15402 17663
rect 15402 17629 15436 17663
rect 15384 17620 15436 17629
rect 15568 17620 15620 17672
rect 11152 17484 11204 17536
rect 14740 17552 14792 17604
rect 14464 17484 14516 17536
rect 14556 17484 14608 17536
rect 3737 17382 3789 17434
rect 3801 17382 3853 17434
rect 3865 17382 3917 17434
rect 3929 17382 3981 17434
rect 3993 17382 4045 17434
rect 7992 17382 8044 17434
rect 8056 17382 8108 17434
rect 8120 17382 8172 17434
rect 8184 17382 8236 17434
rect 8248 17382 8300 17434
rect 12247 17382 12299 17434
rect 12311 17382 12363 17434
rect 12375 17382 12427 17434
rect 12439 17382 12491 17434
rect 12503 17382 12555 17434
rect 16502 17382 16554 17434
rect 16566 17382 16618 17434
rect 16630 17382 16682 17434
rect 16694 17382 16746 17434
rect 16758 17382 16810 17434
rect 4712 17280 4764 17332
rect 5264 17280 5316 17332
rect 4896 17212 4948 17264
rect 2872 17187 2924 17196
rect 2872 17153 2906 17187
rect 2906 17153 2924 17187
rect 2872 17144 2924 17153
rect 6000 17187 6052 17196
rect 6000 17153 6009 17187
rect 6009 17153 6043 17187
rect 6043 17153 6052 17187
rect 6000 17144 6052 17153
rect 9864 17280 9916 17332
rect 10232 17323 10284 17332
rect 10232 17289 10241 17323
rect 10241 17289 10275 17323
rect 10275 17289 10284 17323
rect 10232 17280 10284 17289
rect 14464 17323 14516 17332
rect 14464 17289 14473 17323
rect 14473 17289 14507 17323
rect 14507 17289 14516 17323
rect 14464 17280 14516 17289
rect 14556 17323 14608 17332
rect 14556 17289 14565 17323
rect 14565 17289 14599 17323
rect 14599 17289 14608 17323
rect 14556 17280 14608 17289
rect 15660 17280 15712 17332
rect 7840 17144 7892 17196
rect 8484 17144 8536 17196
rect 2964 16940 3016 16992
rect 5632 17076 5684 17128
rect 7748 17119 7800 17128
rect 7748 17085 7757 17119
rect 7757 17085 7791 17119
rect 7791 17085 7800 17119
rect 7748 17076 7800 17085
rect 8392 17076 8444 17128
rect 10876 17212 10928 17264
rect 15108 17212 15160 17264
rect 11336 17119 11388 17128
rect 11336 17085 11345 17119
rect 11345 17085 11379 17119
rect 11379 17085 11388 17119
rect 11336 17076 11388 17085
rect 13176 17076 13228 17128
rect 5540 16940 5592 16992
rect 10692 16983 10744 16992
rect 10692 16949 10701 16983
rect 10701 16949 10735 16983
rect 10735 16949 10744 16983
rect 10692 16940 10744 16949
rect 3077 16838 3129 16890
rect 3141 16838 3193 16890
rect 3205 16838 3257 16890
rect 3269 16838 3321 16890
rect 3333 16838 3385 16890
rect 7332 16838 7384 16890
rect 7396 16838 7448 16890
rect 7460 16838 7512 16890
rect 7524 16838 7576 16890
rect 7588 16838 7640 16890
rect 11587 16838 11639 16890
rect 11651 16838 11703 16890
rect 11715 16838 11767 16890
rect 11779 16838 11831 16890
rect 11843 16838 11895 16890
rect 15842 16838 15894 16890
rect 15906 16838 15958 16890
rect 15970 16838 16022 16890
rect 16034 16838 16086 16890
rect 16098 16838 16150 16890
rect 2872 16736 2924 16788
rect 5080 16736 5132 16788
rect 2504 16600 2556 16652
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 5172 16643 5224 16652
rect 5172 16609 5181 16643
rect 5181 16609 5215 16643
rect 5215 16609 5224 16643
rect 5172 16600 5224 16609
rect 8668 16736 8720 16788
rect 5540 16600 5592 16652
rect 9588 16600 9640 16652
rect 11060 16736 11112 16788
rect 11336 16736 11388 16788
rect 11980 16600 12032 16652
rect 12532 16643 12584 16652
rect 12532 16609 12541 16643
rect 12541 16609 12575 16643
rect 12575 16609 12584 16643
rect 12532 16600 12584 16609
rect 12900 16643 12952 16652
rect 12900 16609 12934 16643
rect 12934 16609 12952 16643
rect 12900 16600 12952 16609
rect 13084 16643 13136 16652
rect 13084 16609 13093 16643
rect 13093 16609 13127 16643
rect 13127 16609 13136 16643
rect 13084 16600 13136 16609
rect 14464 16600 14516 16652
rect 848 16464 900 16516
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 4252 16575 4304 16584
rect 4252 16541 4261 16575
rect 4261 16541 4295 16575
rect 4295 16541 4304 16575
rect 4252 16532 4304 16541
rect 6920 16575 6972 16584
rect 6920 16541 6929 16575
rect 6929 16541 6963 16575
rect 6963 16541 6972 16575
rect 6920 16532 6972 16541
rect 7748 16532 7800 16584
rect 8760 16532 8812 16584
rect 10232 16532 10284 16584
rect 10876 16532 10928 16584
rect 11612 16532 11664 16584
rect 12072 16575 12124 16584
rect 12072 16541 12081 16575
rect 12081 16541 12115 16575
rect 12115 16541 12124 16575
rect 12072 16532 12124 16541
rect 12808 16575 12860 16584
rect 12808 16541 12817 16575
rect 12817 16541 12851 16575
rect 12851 16541 12860 16575
rect 12808 16532 12860 16541
rect 15292 16575 15344 16584
rect 15292 16541 15301 16575
rect 15301 16541 15335 16575
rect 15335 16541 15344 16575
rect 15292 16532 15344 16541
rect 7196 16507 7248 16516
rect 7196 16473 7230 16507
rect 7230 16473 7248 16507
rect 7196 16464 7248 16473
rect 5448 16396 5500 16448
rect 9220 16464 9272 16516
rect 11520 16464 11572 16516
rect 15568 16643 15620 16652
rect 15568 16609 15577 16643
rect 15577 16609 15611 16643
rect 15611 16609 15620 16643
rect 15568 16600 15620 16609
rect 8944 16439 8996 16448
rect 8944 16405 8953 16439
rect 8953 16405 8987 16439
rect 8987 16405 8996 16439
rect 8944 16396 8996 16405
rect 12072 16396 12124 16448
rect 17040 16439 17092 16448
rect 17040 16405 17049 16439
rect 17049 16405 17083 16439
rect 17083 16405 17092 16439
rect 17040 16396 17092 16405
rect 3737 16294 3789 16346
rect 3801 16294 3853 16346
rect 3865 16294 3917 16346
rect 3929 16294 3981 16346
rect 3993 16294 4045 16346
rect 7992 16294 8044 16346
rect 8056 16294 8108 16346
rect 8120 16294 8172 16346
rect 8184 16294 8236 16346
rect 8248 16294 8300 16346
rect 12247 16294 12299 16346
rect 12311 16294 12363 16346
rect 12375 16294 12427 16346
rect 12439 16294 12491 16346
rect 12503 16294 12555 16346
rect 16502 16294 16554 16346
rect 16566 16294 16618 16346
rect 16630 16294 16682 16346
rect 16694 16294 16746 16346
rect 16758 16294 16810 16346
rect 7196 16235 7248 16244
rect 7196 16201 7205 16235
rect 7205 16201 7239 16235
rect 7239 16201 7248 16235
rect 7196 16192 7248 16201
rect 8944 16192 8996 16244
rect 9220 16192 9272 16244
rect 10600 16192 10652 16244
rect 10692 16192 10744 16244
rect 4436 16124 4488 16176
rect 2964 16056 3016 16108
rect 3424 16099 3476 16108
rect 3424 16065 3458 16099
rect 3458 16065 3476 16099
rect 3424 16056 3476 16065
rect 5356 16056 5408 16108
rect 5816 16056 5868 16108
rect 5264 15920 5316 15972
rect 5724 15920 5776 15972
rect 7840 15988 7892 16040
rect 8760 16124 8812 16176
rect 11152 16124 11204 16176
rect 9588 16099 9640 16108
rect 9588 16065 9622 16099
rect 9622 16065 9640 16099
rect 11520 16235 11572 16244
rect 11520 16201 11529 16235
rect 11529 16201 11563 16235
rect 11563 16201 11572 16235
rect 11520 16192 11572 16201
rect 11612 16192 11664 16244
rect 9588 16056 9640 16065
rect 4620 15895 4672 15904
rect 4620 15861 4629 15895
rect 4629 15861 4663 15895
rect 4663 15861 4672 15895
rect 4620 15852 4672 15861
rect 4712 15852 4764 15904
rect 6092 15852 6144 15904
rect 8944 15988 8996 16040
rect 9312 15988 9364 16040
rect 9496 16031 9548 16040
rect 9496 15997 9505 16031
rect 9505 15997 9539 16031
rect 9539 15997 9548 16031
rect 9496 15988 9548 15997
rect 9956 15988 10008 16040
rect 11888 16099 11940 16108
rect 11888 16065 11897 16099
rect 11897 16065 11931 16099
rect 11931 16065 11940 16099
rect 11888 16056 11940 16065
rect 12072 16099 12124 16108
rect 12072 16065 12081 16099
rect 12081 16065 12115 16099
rect 12115 16065 12124 16099
rect 12072 16056 12124 16065
rect 12808 16099 12860 16108
rect 12808 16065 12817 16099
rect 12817 16065 12851 16099
rect 12851 16065 12860 16099
rect 12808 16056 12860 16065
rect 12900 16099 12952 16108
rect 12900 16065 12934 16099
rect 12934 16065 12952 16099
rect 12900 16056 12952 16065
rect 9220 15963 9272 15972
rect 9220 15929 9229 15963
rect 9229 15929 9263 15963
rect 9263 15929 9272 15963
rect 9220 15920 9272 15929
rect 10232 15920 10284 15972
rect 10692 15920 10744 15972
rect 12532 15963 12584 15972
rect 9128 15852 9180 15904
rect 10140 15852 10192 15904
rect 10324 15852 10376 15904
rect 10600 15852 10652 15904
rect 12532 15929 12541 15963
rect 12541 15929 12575 15963
rect 12575 15929 12584 15963
rect 12532 15920 12584 15929
rect 13268 15852 13320 15904
rect 15292 16192 15344 16244
rect 17040 16192 17092 16244
rect 14924 16124 14976 16176
rect 15200 16056 15252 16108
rect 15660 15920 15712 15972
rect 16488 15988 16540 16040
rect 14740 15852 14792 15904
rect 15752 15852 15804 15904
rect 17684 15895 17736 15904
rect 17684 15861 17693 15895
rect 17693 15861 17727 15895
rect 17727 15861 17736 15895
rect 17684 15852 17736 15861
rect 3077 15750 3129 15802
rect 3141 15750 3193 15802
rect 3205 15750 3257 15802
rect 3269 15750 3321 15802
rect 3333 15750 3385 15802
rect 7332 15750 7384 15802
rect 7396 15750 7448 15802
rect 7460 15750 7512 15802
rect 7524 15750 7576 15802
rect 7588 15750 7640 15802
rect 11587 15750 11639 15802
rect 11651 15750 11703 15802
rect 11715 15750 11767 15802
rect 11779 15750 11831 15802
rect 11843 15750 11895 15802
rect 15842 15750 15894 15802
rect 15906 15750 15958 15802
rect 15970 15750 16022 15802
rect 16034 15750 16086 15802
rect 16098 15750 16150 15802
rect 3424 15691 3476 15700
rect 3424 15657 3433 15691
rect 3433 15657 3467 15691
rect 3467 15657 3476 15691
rect 3424 15648 3476 15657
rect 4712 15648 4764 15700
rect 2504 15512 2556 15564
rect 4252 15555 4304 15564
rect 4252 15521 4261 15555
rect 4261 15521 4295 15555
rect 4295 15521 4304 15555
rect 4252 15512 4304 15521
rect 4436 15555 4488 15564
rect 4436 15521 4445 15555
rect 4445 15521 4479 15555
rect 4479 15521 4488 15555
rect 4436 15512 4488 15521
rect 4620 15444 4672 15496
rect 4712 15444 4764 15496
rect 5540 15648 5592 15700
rect 9496 15648 9548 15700
rect 9864 15648 9916 15700
rect 5448 15555 5500 15564
rect 5448 15521 5457 15555
rect 5457 15521 5491 15555
rect 5491 15521 5500 15555
rect 5448 15512 5500 15521
rect 5816 15555 5868 15564
rect 5816 15521 5850 15555
rect 5850 15521 5868 15555
rect 5816 15512 5868 15521
rect 7104 15512 7156 15564
rect 8944 15555 8996 15564
rect 8944 15521 8953 15555
rect 8953 15521 8987 15555
rect 8987 15521 8996 15555
rect 8944 15512 8996 15521
rect 9128 15555 9180 15564
rect 9128 15521 9137 15555
rect 9137 15521 9171 15555
rect 9171 15521 9180 15555
rect 9128 15512 9180 15521
rect 4896 15444 4948 15496
rect 4252 15376 4304 15428
rect 1492 15351 1544 15360
rect 1492 15317 1501 15351
rect 1501 15317 1535 15351
rect 1535 15317 1544 15351
rect 1492 15308 1544 15317
rect 5172 15444 5224 15496
rect 5724 15487 5776 15496
rect 5724 15453 5733 15487
rect 5733 15453 5767 15487
rect 5767 15453 5776 15487
rect 5724 15444 5776 15453
rect 7656 15444 7708 15496
rect 9680 15512 9732 15564
rect 9864 15487 9916 15496
rect 9864 15453 9873 15487
rect 9873 15453 9907 15487
rect 9907 15453 9916 15487
rect 9864 15444 9916 15453
rect 12532 15512 12584 15564
rect 15568 15512 15620 15564
rect 12716 15444 12768 15496
rect 13084 15444 13136 15496
rect 13912 15444 13964 15496
rect 14740 15487 14792 15496
rect 14740 15453 14749 15487
rect 14749 15453 14783 15487
rect 14783 15453 14792 15487
rect 14740 15444 14792 15453
rect 14832 15444 14884 15496
rect 15016 15487 15068 15496
rect 15016 15453 15025 15487
rect 15025 15453 15059 15487
rect 15059 15453 15068 15487
rect 15016 15444 15068 15453
rect 15844 15444 15896 15496
rect 16120 15444 16172 15496
rect 17500 15487 17552 15496
rect 17500 15453 17509 15487
rect 17509 15453 17543 15487
rect 17543 15453 17552 15487
rect 17500 15444 17552 15453
rect 5632 15308 5684 15360
rect 5724 15308 5776 15360
rect 6644 15351 6696 15360
rect 6644 15317 6653 15351
rect 6653 15317 6687 15351
rect 6687 15317 6696 15351
rect 6644 15308 6696 15317
rect 7288 15351 7340 15360
rect 7288 15317 7297 15351
rect 7297 15317 7331 15351
rect 7331 15317 7340 15351
rect 7288 15308 7340 15317
rect 12808 15376 12860 15428
rect 13728 15376 13780 15428
rect 16304 15419 16356 15428
rect 16304 15385 16338 15419
rect 16338 15385 16356 15419
rect 16304 15376 16356 15385
rect 10784 15351 10836 15360
rect 10784 15317 10793 15351
rect 10793 15317 10827 15351
rect 10827 15317 10836 15351
rect 10784 15308 10836 15317
rect 12624 15308 12676 15360
rect 14280 15308 14332 15360
rect 15844 15308 15896 15360
rect 16488 15308 16540 15360
rect 17684 15351 17736 15360
rect 17684 15317 17693 15351
rect 17693 15317 17727 15351
rect 17727 15317 17736 15351
rect 17684 15308 17736 15317
rect 3737 15206 3789 15258
rect 3801 15206 3853 15258
rect 3865 15206 3917 15258
rect 3929 15206 3981 15258
rect 3993 15206 4045 15258
rect 7992 15206 8044 15258
rect 8056 15206 8108 15258
rect 8120 15206 8172 15258
rect 8184 15206 8236 15258
rect 8248 15206 8300 15258
rect 12247 15206 12299 15258
rect 12311 15206 12363 15258
rect 12375 15206 12427 15258
rect 12439 15206 12491 15258
rect 12503 15206 12555 15258
rect 16502 15206 16554 15258
rect 16566 15206 16618 15258
rect 16630 15206 16682 15258
rect 16694 15206 16746 15258
rect 16758 15206 16810 15258
rect 9772 15104 9824 15156
rect 10508 15147 10560 15156
rect 10508 15113 10517 15147
rect 10517 15113 10551 15147
rect 10551 15113 10560 15147
rect 10508 15104 10560 15113
rect 7288 15036 7340 15088
rect 8668 15036 8720 15088
rect 13912 15104 13964 15156
rect 14832 15104 14884 15156
rect 15752 15104 15804 15156
rect 1768 15011 1820 15020
rect 1768 14977 1802 15011
rect 1802 14977 1820 15011
rect 1768 14968 1820 14977
rect 4712 14968 4764 15020
rect 5264 15011 5316 15020
rect 5264 14977 5273 15011
rect 5273 14977 5307 15011
rect 5307 14977 5316 15011
rect 5264 14968 5316 14977
rect 5356 15011 5408 15020
rect 5356 14977 5390 15011
rect 5390 14977 5408 15011
rect 5356 14968 5408 14977
rect 6552 15011 6604 15020
rect 6552 14977 6561 15011
rect 6561 14977 6595 15011
rect 6595 14977 6604 15011
rect 6552 14968 6604 14977
rect 6644 14968 6696 15020
rect 8484 14968 8536 15020
rect 1400 14900 1452 14952
rect 2780 14832 2832 14884
rect 4896 14900 4948 14952
rect 5724 14900 5776 14952
rect 6920 14943 6972 14952
rect 6920 14909 6929 14943
rect 6929 14909 6963 14943
rect 6963 14909 6972 14943
rect 6920 14900 6972 14909
rect 9312 15011 9364 15020
rect 9312 14977 9321 15011
rect 9321 14977 9355 15011
rect 9355 14977 9364 15011
rect 9312 14968 9364 14977
rect 10232 14968 10284 15020
rect 10324 15011 10376 15020
rect 10324 14977 10333 15011
rect 10333 14977 10367 15011
rect 10367 14977 10376 15011
rect 10324 14968 10376 14977
rect 10508 14968 10560 15020
rect 10784 14968 10836 15020
rect 10968 15011 11020 15020
rect 10968 14977 10977 15011
rect 10977 14977 11011 15011
rect 11011 14977 11020 15011
rect 10968 14968 11020 14977
rect 11152 15011 11204 15020
rect 11152 14977 11161 15011
rect 11161 14977 11195 15011
rect 11195 14977 11204 15011
rect 11152 14968 11204 14977
rect 13912 15011 13964 15020
rect 13912 14977 13930 15011
rect 13930 14977 13964 15011
rect 13912 14968 13964 14977
rect 3516 14764 3568 14816
rect 10048 14832 10100 14884
rect 5448 14764 5500 14816
rect 6184 14807 6236 14816
rect 6184 14773 6193 14807
rect 6193 14773 6227 14807
rect 6227 14773 6236 14807
rect 6184 14764 6236 14773
rect 6368 14807 6420 14816
rect 6368 14773 6377 14807
rect 6377 14773 6411 14807
rect 6411 14773 6420 14807
rect 6368 14764 6420 14773
rect 8392 14807 8444 14816
rect 8392 14773 8401 14807
rect 8401 14773 8435 14807
rect 8435 14773 8444 14807
rect 8392 14764 8444 14773
rect 9220 14764 9272 14816
rect 11060 14900 11112 14952
rect 12716 14900 12768 14952
rect 15016 14968 15068 15020
rect 16120 14968 16172 15020
rect 16304 15147 16356 15156
rect 16304 15113 16313 15147
rect 16313 15113 16347 15147
rect 16347 15113 16356 15147
rect 16304 15104 16356 15113
rect 17776 15011 17828 15020
rect 17776 14977 17785 15011
rect 17785 14977 17819 15011
rect 17819 14977 17828 15011
rect 17776 14968 17828 14977
rect 14372 14832 14424 14884
rect 15660 14943 15712 14952
rect 15660 14909 15669 14943
rect 15669 14909 15703 14943
rect 15703 14909 15712 14943
rect 15660 14900 15712 14909
rect 15844 14832 15896 14884
rect 12164 14764 12216 14816
rect 14740 14764 14792 14816
rect 15108 14764 15160 14816
rect 15660 14764 15712 14816
rect 16396 14900 16448 14952
rect 16856 14807 16908 14816
rect 16856 14773 16865 14807
rect 16865 14773 16899 14807
rect 16899 14773 16908 14807
rect 16856 14764 16908 14773
rect 17592 14807 17644 14816
rect 17592 14773 17601 14807
rect 17601 14773 17635 14807
rect 17635 14773 17644 14807
rect 17592 14764 17644 14773
rect 3077 14662 3129 14714
rect 3141 14662 3193 14714
rect 3205 14662 3257 14714
rect 3269 14662 3321 14714
rect 3333 14662 3385 14714
rect 7332 14662 7384 14714
rect 7396 14662 7448 14714
rect 7460 14662 7512 14714
rect 7524 14662 7576 14714
rect 7588 14662 7640 14714
rect 11587 14662 11639 14714
rect 11651 14662 11703 14714
rect 11715 14662 11767 14714
rect 11779 14662 11831 14714
rect 11843 14662 11895 14714
rect 15842 14662 15894 14714
rect 15906 14662 15958 14714
rect 15970 14662 16022 14714
rect 16034 14662 16086 14714
rect 16098 14662 16150 14714
rect 1768 14560 1820 14612
rect 6092 14603 6144 14612
rect 6092 14569 6101 14603
rect 6101 14569 6135 14603
rect 6135 14569 6144 14603
rect 6092 14560 6144 14569
rect 6184 14560 6236 14612
rect 10140 14560 10192 14612
rect 848 14492 900 14544
rect 6368 14492 6420 14544
rect 10968 14560 11020 14612
rect 2320 14424 2372 14476
rect 8668 14424 8720 14476
rect 11060 14424 11112 14476
rect 11336 14424 11388 14476
rect 2780 14356 2832 14408
rect 6276 14399 6328 14408
rect 6276 14365 6285 14399
rect 6285 14365 6319 14399
rect 6319 14365 6328 14399
rect 6276 14356 6328 14365
rect 6920 14288 6972 14340
rect 9220 14399 9272 14408
rect 9220 14365 9254 14399
rect 9254 14365 9272 14399
rect 9220 14356 9272 14365
rect 14096 14603 14148 14612
rect 14096 14569 14105 14603
rect 14105 14569 14139 14603
rect 14139 14569 14148 14603
rect 14096 14560 14148 14569
rect 14464 14603 14516 14612
rect 14464 14569 14473 14603
rect 14473 14569 14507 14603
rect 14507 14569 14516 14603
rect 14464 14560 14516 14569
rect 14740 14603 14792 14612
rect 14740 14569 14749 14603
rect 14749 14569 14783 14603
rect 14783 14569 14792 14603
rect 14740 14560 14792 14569
rect 15200 14560 15252 14612
rect 17776 14560 17828 14612
rect 16396 14535 16448 14544
rect 16396 14501 16405 14535
rect 16405 14501 16439 14535
rect 16439 14501 16448 14535
rect 16396 14492 16448 14501
rect 15752 14467 15804 14476
rect 15752 14433 15761 14467
rect 15761 14433 15795 14467
rect 15795 14433 15804 14467
rect 15752 14424 15804 14433
rect 13452 14356 13504 14408
rect 14372 14356 14424 14408
rect 8760 14331 8812 14340
rect 8760 14297 8769 14331
rect 8769 14297 8803 14331
rect 8803 14297 8812 14331
rect 8760 14288 8812 14297
rect 13728 14288 13780 14340
rect 15660 14288 15712 14340
rect 16856 14288 16908 14340
rect 17592 14288 17644 14340
rect 2504 14220 2556 14272
rect 8944 14220 8996 14272
rect 12072 14220 12124 14272
rect 15476 14220 15528 14272
rect 16212 14220 16264 14272
rect 3737 14118 3789 14170
rect 3801 14118 3853 14170
rect 3865 14118 3917 14170
rect 3929 14118 3981 14170
rect 3993 14118 4045 14170
rect 7992 14118 8044 14170
rect 8056 14118 8108 14170
rect 8120 14118 8172 14170
rect 8184 14118 8236 14170
rect 8248 14118 8300 14170
rect 12247 14118 12299 14170
rect 12311 14118 12363 14170
rect 12375 14118 12427 14170
rect 12439 14118 12491 14170
rect 12503 14118 12555 14170
rect 16502 14118 16554 14170
rect 16566 14118 16618 14170
rect 16630 14118 16682 14170
rect 16694 14118 16746 14170
rect 16758 14118 16810 14170
rect 6552 14016 6604 14068
rect 7656 14016 7708 14068
rect 8392 14016 8444 14068
rect 2964 13948 3016 14000
rect 4068 13948 4120 14000
rect 4436 13948 4488 14000
rect 1952 13923 2004 13932
rect 1952 13889 1961 13923
rect 1961 13889 1995 13923
rect 1995 13889 2004 13923
rect 1952 13880 2004 13889
rect 5172 13880 5224 13932
rect 6460 13880 6512 13932
rect 3424 13812 3476 13864
rect 6828 13880 6880 13932
rect 7104 13948 7156 14000
rect 8944 13991 8996 14000
rect 8944 13957 8953 13991
rect 8953 13957 8987 13991
rect 8987 13957 8996 13991
rect 8944 13948 8996 13957
rect 7840 13880 7892 13932
rect 7932 13923 7984 13932
rect 7932 13889 7941 13923
rect 7941 13889 7975 13923
rect 7975 13889 7984 13923
rect 9312 14059 9364 14068
rect 9312 14025 9321 14059
rect 9321 14025 9355 14059
rect 9355 14025 9364 14059
rect 9312 14016 9364 14025
rect 10048 14059 10100 14068
rect 10048 14025 10057 14059
rect 10057 14025 10091 14059
rect 10091 14025 10100 14059
rect 10048 14016 10100 14025
rect 10140 14059 10192 14068
rect 10140 14025 10149 14059
rect 10149 14025 10183 14059
rect 10183 14025 10192 14059
rect 10140 14016 10192 14025
rect 11152 14016 11204 14068
rect 12624 14016 12676 14068
rect 13544 14016 13596 14068
rect 16396 14016 16448 14068
rect 16948 14059 17000 14068
rect 16948 14025 16957 14059
rect 16957 14025 16991 14059
rect 16991 14025 17000 14059
rect 16948 14016 17000 14025
rect 12072 13991 12124 14000
rect 12072 13957 12081 13991
rect 12081 13957 12115 13991
rect 12115 13957 12124 13991
rect 12072 13948 12124 13957
rect 12164 13948 12216 14000
rect 7932 13880 7984 13889
rect 9956 13880 10008 13932
rect 12624 13923 12676 13932
rect 12624 13889 12633 13923
rect 12633 13889 12667 13923
rect 12667 13889 12676 13923
rect 12624 13880 12676 13889
rect 13268 13923 13320 13932
rect 13268 13889 13277 13923
rect 13277 13889 13311 13923
rect 13311 13889 13320 13923
rect 13268 13880 13320 13889
rect 13912 13880 13964 13932
rect 14280 13923 14332 13932
rect 14280 13889 14289 13923
rect 14289 13889 14323 13923
rect 14323 13889 14332 13923
rect 14280 13880 14332 13889
rect 14464 13923 14516 13932
rect 14464 13889 14473 13923
rect 14473 13889 14507 13923
rect 14507 13889 14516 13923
rect 14464 13880 14516 13889
rect 2964 13744 3016 13796
rect 1676 13676 1728 13728
rect 2688 13719 2740 13728
rect 2688 13685 2697 13719
rect 2697 13685 2731 13719
rect 2731 13685 2740 13719
rect 2688 13676 2740 13685
rect 5540 13719 5592 13728
rect 5540 13685 5549 13719
rect 5549 13685 5583 13719
rect 5583 13685 5592 13719
rect 5540 13676 5592 13685
rect 7656 13744 7708 13796
rect 8576 13744 8628 13796
rect 9864 13812 9916 13864
rect 10692 13812 10744 13864
rect 11152 13812 11204 13864
rect 9680 13719 9732 13728
rect 9680 13685 9689 13719
rect 9689 13685 9723 13719
rect 9723 13685 9732 13719
rect 9680 13676 9732 13685
rect 12440 13719 12492 13728
rect 12440 13685 12449 13719
rect 12449 13685 12483 13719
rect 12483 13685 12492 13719
rect 12440 13676 12492 13685
rect 15292 13948 15344 14000
rect 16304 13948 16356 14000
rect 15200 13855 15252 13864
rect 15200 13821 15209 13855
rect 15209 13821 15243 13855
rect 15243 13821 15252 13855
rect 15200 13812 15252 13821
rect 15108 13744 15160 13796
rect 15660 13812 15712 13864
rect 14556 13676 14608 13728
rect 14648 13719 14700 13728
rect 14648 13685 14657 13719
rect 14657 13685 14691 13719
rect 14691 13685 14700 13719
rect 14648 13676 14700 13685
rect 15200 13676 15252 13728
rect 17132 13719 17184 13728
rect 17132 13685 17141 13719
rect 17141 13685 17175 13719
rect 17175 13685 17184 13719
rect 17132 13676 17184 13685
rect 3077 13574 3129 13626
rect 3141 13574 3193 13626
rect 3205 13574 3257 13626
rect 3269 13574 3321 13626
rect 3333 13574 3385 13626
rect 7332 13574 7384 13626
rect 7396 13574 7448 13626
rect 7460 13574 7512 13626
rect 7524 13574 7576 13626
rect 7588 13574 7640 13626
rect 11587 13574 11639 13626
rect 11651 13574 11703 13626
rect 11715 13574 11767 13626
rect 11779 13574 11831 13626
rect 11843 13574 11895 13626
rect 15842 13574 15894 13626
rect 15906 13574 15958 13626
rect 15970 13574 16022 13626
rect 16034 13574 16086 13626
rect 16098 13574 16150 13626
rect 3056 13472 3108 13524
rect 3056 13379 3108 13388
rect 3056 13345 3065 13379
rect 3065 13345 3099 13379
rect 3099 13345 3108 13379
rect 3056 13336 3108 13345
rect 3424 13336 3476 13388
rect 4068 13336 4120 13388
rect 10508 13472 10560 13524
rect 15568 13472 15620 13524
rect 16212 13472 16264 13524
rect 5724 13404 5776 13456
rect 10140 13404 10192 13456
rect 10232 13336 10284 13388
rect 1400 13311 1452 13320
rect 1400 13277 1409 13311
rect 1409 13277 1443 13311
rect 1443 13277 1452 13311
rect 1400 13268 1452 13277
rect 1676 13311 1728 13320
rect 1676 13277 1710 13311
rect 1710 13277 1728 13311
rect 1676 13268 1728 13277
rect 2780 13268 2832 13320
rect 3516 13268 3568 13320
rect 6000 13311 6052 13320
rect 6000 13277 6009 13311
rect 6009 13277 6043 13311
rect 6043 13277 6052 13311
rect 6000 13268 6052 13277
rect 6552 13311 6604 13320
rect 6552 13277 6561 13311
rect 6561 13277 6595 13311
rect 6595 13277 6604 13311
rect 6552 13268 6604 13277
rect 6736 13268 6788 13320
rect 7104 13268 7156 13320
rect 10324 13268 10376 13320
rect 10600 13311 10652 13320
rect 10600 13277 10604 13311
rect 10604 13277 10638 13311
rect 10638 13277 10652 13311
rect 10600 13268 10652 13277
rect 10692 13311 10744 13320
rect 10692 13277 10701 13311
rect 10701 13277 10735 13311
rect 10735 13277 10744 13311
rect 10692 13268 10744 13277
rect 2596 13200 2648 13252
rect 8576 13200 8628 13252
rect 10048 13200 10100 13252
rect 10140 13200 10192 13252
rect 11336 13379 11388 13388
rect 11336 13345 11345 13379
rect 11345 13345 11379 13379
rect 11379 13345 11388 13379
rect 11336 13336 11388 13345
rect 14648 13404 14700 13456
rect 17500 13404 17552 13456
rect 12992 13336 13044 13388
rect 17224 13336 17276 13388
rect 12440 13268 12492 13320
rect 13820 13268 13872 13320
rect 15476 13268 15528 13320
rect 5816 13132 5868 13184
rect 6368 13175 6420 13184
rect 6368 13141 6377 13175
rect 6377 13141 6411 13175
rect 6411 13141 6420 13175
rect 6368 13132 6420 13141
rect 6644 13132 6696 13184
rect 8944 13132 8996 13184
rect 13268 13200 13320 13252
rect 13360 13200 13412 13252
rect 15568 13200 15620 13252
rect 17132 13268 17184 13320
rect 17684 13243 17736 13252
rect 17684 13209 17693 13243
rect 17693 13209 17727 13243
rect 17727 13209 17736 13243
rect 17684 13200 17736 13209
rect 12808 13175 12860 13184
rect 12808 13141 12817 13175
rect 12817 13141 12851 13175
rect 12851 13141 12860 13175
rect 12808 13132 12860 13141
rect 14648 13132 14700 13184
rect 15660 13132 15712 13184
rect 17500 13132 17552 13184
rect 3737 13030 3789 13082
rect 3801 13030 3853 13082
rect 3865 13030 3917 13082
rect 3929 13030 3981 13082
rect 3993 13030 4045 13082
rect 7992 13030 8044 13082
rect 8056 13030 8108 13082
rect 8120 13030 8172 13082
rect 8184 13030 8236 13082
rect 8248 13030 8300 13082
rect 12247 13030 12299 13082
rect 12311 13030 12363 13082
rect 12375 13030 12427 13082
rect 12439 13030 12491 13082
rect 12503 13030 12555 13082
rect 16502 13030 16554 13082
rect 16566 13030 16618 13082
rect 16630 13030 16682 13082
rect 16694 13030 16746 13082
rect 16758 13030 16810 13082
rect 1952 12928 2004 12980
rect 2688 12928 2740 12980
rect 3424 12928 3476 12980
rect 1032 12860 1084 12912
rect 3516 12860 3568 12912
rect 2504 12724 2556 12776
rect 2688 12767 2740 12776
rect 2688 12733 2697 12767
rect 2697 12733 2731 12767
rect 2731 12733 2740 12767
rect 2688 12724 2740 12733
rect 2964 12724 3016 12776
rect 1400 12656 1452 12708
rect 2872 12656 2924 12708
rect 3700 12792 3752 12844
rect 3884 12792 3936 12844
rect 4068 12835 4120 12844
rect 4068 12801 4102 12835
rect 4102 12801 4120 12835
rect 4068 12792 4120 12801
rect 5540 12928 5592 12980
rect 6276 12928 6328 12980
rect 5816 12903 5868 12912
rect 5816 12869 5825 12903
rect 5825 12869 5859 12903
rect 5859 12869 5868 12903
rect 5816 12860 5868 12869
rect 9680 12860 9732 12912
rect 10416 12971 10468 12980
rect 10416 12937 10425 12971
rect 10425 12937 10459 12971
rect 10459 12937 10468 12971
rect 10416 12928 10468 12937
rect 12072 12928 12124 12980
rect 12624 12971 12676 12980
rect 12624 12937 12633 12971
rect 12633 12937 12667 12971
rect 12667 12937 12676 12971
rect 12624 12928 12676 12937
rect 14372 12928 14424 12980
rect 14464 12928 14516 12980
rect 5724 12835 5776 12844
rect 5724 12801 5731 12835
rect 5731 12801 5776 12835
rect 5724 12792 5776 12801
rect 5908 12835 5960 12844
rect 5908 12801 5917 12835
rect 5917 12801 5951 12835
rect 5951 12801 5960 12835
rect 5908 12792 5960 12801
rect 6368 12792 6420 12844
rect 7012 12792 7064 12844
rect 9220 12835 9272 12844
rect 9220 12801 9229 12835
rect 9229 12801 9263 12835
rect 9263 12801 9272 12835
rect 9220 12792 9272 12801
rect 6920 12767 6972 12776
rect 6920 12733 6929 12767
rect 6929 12733 6963 12767
rect 6963 12733 6972 12767
rect 6920 12724 6972 12733
rect 5632 12656 5684 12708
rect 6644 12656 6696 12708
rect 4436 12588 4488 12640
rect 7104 12588 7156 12640
rect 9956 12835 10008 12844
rect 9956 12801 9963 12835
rect 9963 12801 10008 12835
rect 9956 12792 10008 12801
rect 10876 12835 10928 12844
rect 10876 12801 10885 12835
rect 10885 12801 10919 12835
rect 10919 12801 10928 12835
rect 10876 12792 10928 12801
rect 11244 12792 11296 12844
rect 12808 12860 12860 12912
rect 13544 12903 13596 12912
rect 13544 12869 13553 12903
rect 13553 12869 13587 12903
rect 13587 12869 13596 12903
rect 13544 12860 13596 12869
rect 15200 12860 15252 12912
rect 12440 12792 12492 12844
rect 12716 12835 12768 12844
rect 12716 12801 12725 12835
rect 12725 12801 12759 12835
rect 12759 12801 12768 12835
rect 12716 12792 12768 12801
rect 13268 12835 13320 12844
rect 13268 12801 13277 12835
rect 13277 12801 13311 12835
rect 13311 12801 13320 12835
rect 13268 12792 13320 12801
rect 13360 12835 13412 12844
rect 13360 12801 13370 12835
rect 13370 12801 13404 12835
rect 13404 12801 13412 12835
rect 13360 12792 13412 12801
rect 12072 12767 12124 12776
rect 12072 12733 12081 12767
rect 12081 12733 12115 12767
rect 12115 12733 12124 12767
rect 12072 12724 12124 12733
rect 13728 12835 13780 12844
rect 13728 12801 13742 12835
rect 13742 12801 13776 12835
rect 13776 12801 13780 12835
rect 13728 12792 13780 12801
rect 14188 12835 14240 12844
rect 14188 12801 14195 12835
rect 14195 12801 14240 12835
rect 14188 12792 14240 12801
rect 14372 12835 14424 12844
rect 14372 12801 14381 12835
rect 14381 12801 14415 12835
rect 14415 12801 14424 12835
rect 14372 12792 14424 12801
rect 14464 12835 14516 12844
rect 14464 12801 14478 12835
rect 14478 12801 14512 12835
rect 14512 12801 14516 12835
rect 14464 12792 14516 12801
rect 16580 12792 16632 12844
rect 14556 12724 14608 12776
rect 16488 12767 16540 12776
rect 16488 12733 16497 12767
rect 16497 12733 16531 12767
rect 16531 12733 16540 12767
rect 16488 12724 16540 12733
rect 8392 12631 8444 12640
rect 8392 12597 8401 12631
rect 8401 12597 8435 12631
rect 8435 12597 8444 12631
rect 8392 12588 8444 12597
rect 9404 12631 9456 12640
rect 9404 12597 9413 12631
rect 9413 12597 9447 12631
rect 9447 12597 9456 12631
rect 9404 12588 9456 12597
rect 9680 12588 9732 12640
rect 10232 12588 10284 12640
rect 12624 12588 12676 12640
rect 12992 12631 13044 12640
rect 12992 12597 13001 12631
rect 13001 12597 13035 12631
rect 13035 12597 13044 12631
rect 12992 12588 13044 12597
rect 14924 12588 14976 12640
rect 16672 12631 16724 12640
rect 16672 12597 16681 12631
rect 16681 12597 16715 12631
rect 16715 12597 16724 12631
rect 16672 12588 16724 12597
rect 3077 12486 3129 12538
rect 3141 12486 3193 12538
rect 3205 12486 3257 12538
rect 3269 12486 3321 12538
rect 3333 12486 3385 12538
rect 7332 12486 7384 12538
rect 7396 12486 7448 12538
rect 7460 12486 7512 12538
rect 7524 12486 7576 12538
rect 7588 12486 7640 12538
rect 11587 12486 11639 12538
rect 11651 12486 11703 12538
rect 11715 12486 11767 12538
rect 11779 12486 11831 12538
rect 11843 12486 11895 12538
rect 15842 12486 15894 12538
rect 15906 12486 15958 12538
rect 15970 12486 16022 12538
rect 16034 12486 16086 12538
rect 16098 12486 16150 12538
rect 4068 12384 4120 12436
rect 5908 12384 5960 12436
rect 2504 12248 2556 12300
rect 1308 12180 1360 12232
rect 2044 12180 2096 12232
rect 2872 12180 2924 12232
rect 1768 12087 1820 12096
rect 1768 12053 1777 12087
rect 1777 12053 1811 12087
rect 1811 12053 1820 12087
rect 1768 12044 1820 12053
rect 1860 12044 1912 12096
rect 2412 12044 2464 12096
rect 4804 12291 4856 12300
rect 4804 12257 4813 12291
rect 4813 12257 4847 12291
rect 4847 12257 4856 12291
rect 4804 12248 4856 12257
rect 5540 12248 5592 12300
rect 6460 12384 6512 12436
rect 7012 12384 7064 12436
rect 6092 12316 6144 12368
rect 7840 12384 7892 12436
rect 8208 12384 8260 12436
rect 6736 12248 6788 12300
rect 8392 12316 8444 12368
rect 9404 12384 9456 12436
rect 10600 12384 10652 12436
rect 12992 12427 13044 12436
rect 12992 12393 13001 12427
rect 13001 12393 13035 12427
rect 13035 12393 13044 12427
rect 12992 12384 13044 12393
rect 13728 12384 13780 12436
rect 16304 12427 16356 12436
rect 16304 12393 16313 12427
rect 16313 12393 16347 12427
rect 16347 12393 16356 12427
rect 16304 12384 16356 12393
rect 16396 12427 16448 12436
rect 16396 12393 16405 12427
rect 16405 12393 16439 12427
rect 16439 12393 16448 12427
rect 16396 12384 16448 12393
rect 9680 12316 9732 12368
rect 14372 12316 14424 12368
rect 5172 12180 5224 12232
rect 5448 12180 5500 12232
rect 6552 12223 6604 12232
rect 6552 12189 6561 12223
rect 6561 12189 6595 12223
rect 6595 12189 6604 12223
rect 6552 12180 6604 12189
rect 7104 12180 7156 12232
rect 7840 12248 7892 12300
rect 8392 12223 8444 12232
rect 8392 12189 8401 12223
rect 8401 12189 8435 12223
rect 8435 12189 8444 12223
rect 8392 12180 8444 12189
rect 8944 12223 8996 12232
rect 8944 12189 8953 12223
rect 8953 12189 8987 12223
rect 8987 12189 8996 12223
rect 8944 12180 8996 12189
rect 10692 12248 10744 12300
rect 15108 12248 15160 12300
rect 15200 12248 15252 12300
rect 16672 12248 16724 12300
rect 7196 12112 7248 12164
rect 9220 12112 9272 12164
rect 11244 12180 11296 12232
rect 12440 12180 12492 12232
rect 12808 12223 12860 12232
rect 12808 12189 12817 12223
rect 12817 12189 12851 12223
rect 12851 12189 12860 12223
rect 12808 12180 12860 12189
rect 13820 12180 13872 12232
rect 12716 12112 12768 12164
rect 8576 12044 8628 12096
rect 9036 12087 9088 12096
rect 9036 12053 9045 12087
rect 9045 12053 9079 12087
rect 9079 12053 9088 12087
rect 9036 12044 9088 12053
rect 12624 12044 12676 12096
rect 14004 12044 14056 12096
rect 14832 12180 14884 12232
rect 14924 12223 14976 12232
rect 14924 12189 14933 12223
rect 14933 12189 14967 12223
rect 14967 12189 14976 12223
rect 14924 12180 14976 12189
rect 16396 12180 16448 12232
rect 15660 12112 15712 12164
rect 17684 12112 17736 12164
rect 3737 11942 3789 11994
rect 3801 11942 3853 11994
rect 3865 11942 3917 11994
rect 3929 11942 3981 11994
rect 3993 11942 4045 11994
rect 7992 11942 8044 11994
rect 8056 11942 8108 11994
rect 8120 11942 8172 11994
rect 8184 11942 8236 11994
rect 8248 11942 8300 11994
rect 12247 11942 12299 11994
rect 12311 11942 12363 11994
rect 12375 11942 12427 11994
rect 12439 11942 12491 11994
rect 12503 11942 12555 11994
rect 16502 11942 16554 11994
rect 16566 11942 16618 11994
rect 16630 11942 16682 11994
rect 16694 11942 16746 11994
rect 16758 11942 16810 11994
rect 4804 11840 4856 11892
rect 8668 11840 8720 11892
rect 1768 11772 1820 11824
rect 5540 11772 5592 11824
rect 1860 11747 1912 11756
rect 1860 11713 1894 11747
rect 1894 11713 1912 11747
rect 1860 11704 1912 11713
rect 3608 11747 3660 11756
rect 3608 11713 3617 11747
rect 3617 11713 3651 11747
rect 3651 11713 3660 11747
rect 3608 11704 3660 11713
rect 3884 11747 3936 11756
rect 3884 11713 3918 11747
rect 3918 11713 3936 11747
rect 3884 11704 3936 11713
rect 6644 11704 6696 11756
rect 6736 11704 6788 11756
rect 7012 11747 7064 11756
rect 7012 11713 7021 11747
rect 7021 11713 7055 11747
rect 7055 11713 7064 11747
rect 7012 11704 7064 11713
rect 9864 11772 9916 11824
rect 10324 11772 10376 11824
rect 11428 11704 11480 11756
rect 12808 11704 12860 11756
rect 13728 11704 13780 11756
rect 14004 11840 14056 11892
rect 14464 11840 14516 11892
rect 17684 11883 17736 11892
rect 17684 11849 17693 11883
rect 17693 11849 17727 11883
rect 17727 11849 17736 11883
rect 17684 11840 17736 11849
rect 14004 11747 14056 11756
rect 14004 11713 14013 11747
rect 14013 11713 14047 11747
rect 14047 11713 14056 11747
rect 14004 11704 14056 11713
rect 14924 11772 14976 11824
rect 15752 11772 15804 11824
rect 1400 11636 1452 11688
rect 5356 11636 5408 11688
rect 4620 11568 4672 11620
rect 5908 11568 5960 11620
rect 6828 11568 6880 11620
rect 8668 11568 8720 11620
rect 9404 11636 9456 11688
rect 14648 11704 14700 11756
rect 15016 11704 15068 11756
rect 2872 11500 2924 11552
rect 5356 11500 5408 11552
rect 6368 11543 6420 11552
rect 6368 11509 6377 11543
rect 6377 11509 6411 11543
rect 6411 11509 6420 11543
rect 6368 11500 6420 11509
rect 8484 11543 8536 11552
rect 8484 11509 8493 11543
rect 8493 11509 8527 11543
rect 8527 11509 8536 11543
rect 8484 11500 8536 11509
rect 13084 11611 13136 11620
rect 13084 11577 13093 11611
rect 13093 11577 13127 11611
rect 13127 11577 13136 11611
rect 13084 11568 13136 11577
rect 13728 11568 13780 11620
rect 17500 11747 17552 11756
rect 17500 11713 17509 11747
rect 17509 11713 17543 11747
rect 17543 11713 17552 11747
rect 17500 11704 17552 11713
rect 16212 11636 16264 11688
rect 17132 11679 17184 11688
rect 17132 11645 17141 11679
rect 17141 11645 17175 11679
rect 17175 11645 17184 11679
rect 17132 11636 17184 11645
rect 17224 11679 17276 11688
rect 17224 11645 17233 11679
rect 17233 11645 17267 11679
rect 17267 11645 17276 11679
rect 17224 11636 17276 11645
rect 11152 11500 11204 11552
rect 12256 11500 12308 11552
rect 12624 11500 12676 11552
rect 13544 11500 13596 11552
rect 15752 11543 15804 11552
rect 15752 11509 15761 11543
rect 15761 11509 15795 11543
rect 15795 11509 15804 11543
rect 15752 11500 15804 11509
rect 3077 11398 3129 11450
rect 3141 11398 3193 11450
rect 3205 11398 3257 11450
rect 3269 11398 3321 11450
rect 3333 11398 3385 11450
rect 7332 11398 7384 11450
rect 7396 11398 7448 11450
rect 7460 11398 7512 11450
rect 7524 11398 7576 11450
rect 7588 11398 7640 11450
rect 11587 11398 11639 11450
rect 11651 11398 11703 11450
rect 11715 11398 11767 11450
rect 11779 11398 11831 11450
rect 11843 11398 11895 11450
rect 15842 11398 15894 11450
rect 15906 11398 15958 11450
rect 15970 11398 16022 11450
rect 16034 11398 16086 11450
rect 16098 11398 16150 11450
rect 2044 11339 2096 11348
rect 2044 11305 2053 11339
rect 2053 11305 2087 11339
rect 2087 11305 2096 11339
rect 2044 11296 2096 11305
rect 3884 11296 3936 11348
rect 5356 11339 5408 11348
rect 5356 11305 5365 11339
rect 5365 11305 5399 11339
rect 5399 11305 5408 11339
rect 5356 11296 5408 11305
rect 6552 11296 6604 11348
rect 2320 11160 2372 11212
rect 1952 11135 2004 11144
rect 1952 11101 1961 11135
rect 1961 11101 1995 11135
rect 1995 11101 2004 11135
rect 1952 11092 2004 11101
rect 2412 11135 2464 11144
rect 2412 11101 2421 11135
rect 2421 11101 2455 11135
rect 2455 11101 2464 11135
rect 2412 11092 2464 11101
rect 2964 11203 3016 11212
rect 2964 11169 2973 11203
rect 2973 11169 3007 11203
rect 3007 11169 3016 11203
rect 2964 11160 3016 11169
rect 3056 11092 3108 11144
rect 5540 11228 5592 11280
rect 6092 11228 6144 11280
rect 4804 11203 4856 11212
rect 4804 11169 4813 11203
rect 4813 11169 4847 11203
rect 4847 11169 4856 11203
rect 4804 11160 4856 11169
rect 4620 11135 4672 11144
rect 4620 11101 4629 11135
rect 4629 11101 4663 11135
rect 4663 11101 4672 11135
rect 4620 11092 4672 11101
rect 4712 11135 4764 11144
rect 4712 11101 4721 11135
rect 4721 11101 4755 11135
rect 4755 11101 4764 11135
rect 4712 11092 4764 11101
rect 5080 11135 5132 11144
rect 5080 11101 5089 11135
rect 5089 11101 5123 11135
rect 5123 11101 5132 11135
rect 5080 11092 5132 11101
rect 5540 11092 5592 11144
rect 5816 11135 5868 11144
rect 5816 11101 5823 11135
rect 5823 11101 5868 11135
rect 5816 11092 5868 11101
rect 1492 11067 1544 11076
rect 1492 11033 1501 11067
rect 1501 11033 1535 11067
rect 1535 11033 1544 11067
rect 1492 11024 1544 11033
rect 1768 10999 1820 11008
rect 1768 10965 1777 10999
rect 1777 10965 1811 10999
rect 1811 10965 1820 10999
rect 1768 10956 1820 10965
rect 2872 11024 2924 11076
rect 2688 10956 2740 11008
rect 3148 10999 3200 11008
rect 3148 10965 3157 10999
rect 3157 10965 3191 10999
rect 3191 10965 3200 10999
rect 3148 10956 3200 10965
rect 3240 10999 3292 11008
rect 3240 10965 3249 10999
rect 3249 10965 3283 10999
rect 3283 10965 3292 10999
rect 3240 10956 3292 10965
rect 6000 11067 6052 11076
rect 6000 11033 6009 11067
rect 6009 11033 6043 11067
rect 6043 11033 6052 11067
rect 6000 11024 6052 11033
rect 9772 11296 9824 11348
rect 13084 11296 13136 11348
rect 14096 11296 14148 11348
rect 12808 11228 12860 11280
rect 14372 11228 14424 11280
rect 14924 11228 14976 11280
rect 7012 11092 7064 11144
rect 7196 11092 7248 11144
rect 7840 11203 7892 11212
rect 7840 11169 7849 11203
rect 7849 11169 7883 11203
rect 7883 11169 7892 11203
rect 7840 11160 7892 11169
rect 15016 11160 15068 11212
rect 16212 11228 16264 11280
rect 9680 11092 9732 11144
rect 11336 11092 11388 11144
rect 12256 11092 12308 11144
rect 12624 11092 12676 11144
rect 16396 11092 16448 11144
rect 5540 10999 5592 11008
rect 5540 10965 5549 10999
rect 5549 10965 5583 10999
rect 5583 10965 5592 10999
rect 5540 10956 5592 10965
rect 6276 10999 6328 11008
rect 6276 10965 6285 10999
rect 6285 10965 6319 10999
rect 6319 10965 6328 10999
rect 6276 10956 6328 10965
rect 7104 10956 7156 11008
rect 7196 10956 7248 11008
rect 12072 11024 12124 11076
rect 11336 10956 11388 11008
rect 12624 10999 12676 11008
rect 12624 10965 12633 10999
rect 12633 10965 12667 10999
rect 12667 10965 12676 10999
rect 12624 10956 12676 10965
rect 14188 10956 14240 11008
rect 15108 10956 15160 11008
rect 15568 10999 15620 11008
rect 15568 10965 15577 10999
rect 15577 10965 15611 10999
rect 15611 10965 15620 10999
rect 15568 10956 15620 10965
rect 15752 11024 15804 11076
rect 16856 10956 16908 11008
rect 3737 10854 3789 10906
rect 3801 10854 3853 10906
rect 3865 10854 3917 10906
rect 3929 10854 3981 10906
rect 3993 10854 4045 10906
rect 7992 10854 8044 10906
rect 8056 10854 8108 10906
rect 8120 10854 8172 10906
rect 8184 10854 8236 10906
rect 8248 10854 8300 10906
rect 12247 10854 12299 10906
rect 12311 10854 12363 10906
rect 12375 10854 12427 10906
rect 12439 10854 12491 10906
rect 12503 10854 12555 10906
rect 16502 10854 16554 10906
rect 16566 10854 16618 10906
rect 16630 10854 16682 10906
rect 16694 10854 16746 10906
rect 16758 10854 16810 10906
rect 3148 10752 3200 10804
rect 3240 10752 3292 10804
rect 1768 10684 1820 10736
rect 5540 10752 5592 10804
rect 7012 10752 7064 10804
rect 9404 10795 9456 10804
rect 9404 10761 9413 10795
rect 9413 10761 9447 10795
rect 9447 10761 9456 10795
rect 9404 10752 9456 10761
rect 10784 10795 10836 10804
rect 10784 10761 10793 10795
rect 10793 10761 10827 10795
rect 10827 10761 10836 10795
rect 10784 10752 10836 10761
rect 11428 10752 11480 10804
rect 12072 10795 12124 10804
rect 12072 10761 12081 10795
rect 12081 10761 12115 10795
rect 12115 10761 12124 10795
rect 12072 10752 12124 10761
rect 13268 10752 13320 10804
rect 13452 10752 13504 10804
rect 13912 10752 13964 10804
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 3148 10616 3200 10668
rect 5264 10616 5316 10668
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 5724 10659 5776 10668
rect 5724 10625 5731 10659
rect 5731 10625 5776 10659
rect 5724 10616 5776 10625
rect 6368 10616 6420 10668
rect 6920 10684 6972 10736
rect 6828 10659 6880 10668
rect 6828 10625 6862 10659
rect 6862 10625 6880 10659
rect 6828 10616 6880 10625
rect 8484 10684 8536 10736
rect 10968 10684 11020 10736
rect 9496 10659 9548 10668
rect 9496 10625 9505 10659
rect 9505 10625 9539 10659
rect 9539 10625 9548 10659
rect 9496 10616 9548 10625
rect 11152 10616 11204 10668
rect 11980 10616 12032 10668
rect 12716 10616 12768 10668
rect 2780 10548 2832 10600
rect 3424 10591 3476 10600
rect 3424 10557 3433 10591
rect 3433 10557 3467 10591
rect 3467 10557 3476 10591
rect 3424 10548 3476 10557
rect 12256 10591 12308 10600
rect 12256 10557 12265 10591
rect 12265 10557 12299 10591
rect 12299 10557 12308 10591
rect 12256 10548 12308 10557
rect 6000 10480 6052 10532
rect 15568 10752 15620 10804
rect 14096 10727 14148 10736
rect 14096 10693 14105 10727
rect 14105 10693 14139 10727
rect 14139 10693 14148 10727
rect 14096 10684 14148 10693
rect 14188 10727 14240 10736
rect 14188 10693 14197 10727
rect 14197 10693 14231 10727
rect 14231 10693 14240 10727
rect 14188 10684 14240 10693
rect 13084 10659 13136 10668
rect 13084 10625 13093 10659
rect 13093 10625 13127 10659
rect 13127 10625 13136 10659
rect 13084 10616 13136 10625
rect 13268 10659 13320 10668
rect 13268 10625 13275 10659
rect 13275 10625 13320 10659
rect 13268 10616 13320 10625
rect 13544 10659 13596 10668
rect 13544 10625 13558 10659
rect 13558 10625 13592 10659
rect 13592 10625 13596 10659
rect 13544 10616 13596 10625
rect 13912 10616 13964 10668
rect 14280 10659 14332 10668
rect 14280 10625 14325 10659
rect 14325 10625 14332 10659
rect 14280 10616 14332 10625
rect 14556 10616 14608 10668
rect 14832 10616 14884 10668
rect 16212 10659 16264 10668
rect 16212 10625 16230 10659
rect 16230 10625 16264 10659
rect 16212 10616 16264 10625
rect 16396 10616 16448 10668
rect 17500 10616 17552 10668
rect 17684 10659 17736 10668
rect 17684 10625 17693 10659
rect 17693 10625 17727 10659
rect 17727 10625 17736 10659
rect 17684 10616 17736 10625
rect 17132 10591 17184 10600
rect 14464 10480 14516 10532
rect 4160 10455 4212 10464
rect 4160 10421 4169 10455
rect 4169 10421 4203 10455
rect 4203 10421 4212 10455
rect 4160 10412 4212 10421
rect 5356 10412 5408 10464
rect 7840 10412 7892 10464
rect 12624 10455 12676 10464
rect 12624 10421 12633 10455
rect 12633 10421 12667 10455
rect 12667 10421 12676 10455
rect 12624 10412 12676 10421
rect 14556 10455 14608 10464
rect 14556 10421 14565 10455
rect 14565 10421 14599 10455
rect 14599 10421 14608 10455
rect 14556 10412 14608 10421
rect 15108 10523 15160 10532
rect 15108 10489 15117 10523
rect 15117 10489 15151 10523
rect 15151 10489 15160 10523
rect 15108 10480 15160 10489
rect 17132 10557 17141 10591
rect 17141 10557 17175 10591
rect 17175 10557 17184 10591
rect 17132 10548 17184 10557
rect 17316 10591 17368 10600
rect 17316 10557 17325 10591
rect 17325 10557 17359 10591
rect 17359 10557 17368 10591
rect 17316 10548 17368 10557
rect 16672 10455 16724 10464
rect 16672 10421 16681 10455
rect 16681 10421 16715 10455
rect 16715 10421 16724 10455
rect 16672 10412 16724 10421
rect 3077 10310 3129 10362
rect 3141 10310 3193 10362
rect 3205 10310 3257 10362
rect 3269 10310 3321 10362
rect 3333 10310 3385 10362
rect 7332 10310 7384 10362
rect 7396 10310 7448 10362
rect 7460 10310 7512 10362
rect 7524 10310 7576 10362
rect 7588 10310 7640 10362
rect 11587 10310 11639 10362
rect 11651 10310 11703 10362
rect 11715 10310 11767 10362
rect 11779 10310 11831 10362
rect 11843 10310 11895 10362
rect 15842 10310 15894 10362
rect 15906 10310 15958 10362
rect 15970 10310 16022 10362
rect 16034 10310 16086 10362
rect 16098 10310 16150 10362
rect 1216 10208 1268 10260
rect 1952 10208 2004 10260
rect 6828 10208 6880 10260
rect 9680 10208 9732 10260
rect 2596 10140 2648 10192
rect 9772 10140 9824 10192
rect 12624 10208 12676 10260
rect 12808 10251 12860 10260
rect 12808 10217 12817 10251
rect 12817 10217 12851 10251
rect 12851 10217 12860 10251
rect 12808 10208 12860 10217
rect 13912 10251 13964 10260
rect 13912 10217 13921 10251
rect 13921 10217 13955 10251
rect 13955 10217 13964 10251
rect 13912 10208 13964 10217
rect 14832 10251 14884 10260
rect 14832 10217 14841 10251
rect 14841 10217 14875 10251
rect 14875 10217 14884 10251
rect 14832 10208 14884 10217
rect 16212 10208 16264 10260
rect 17500 10251 17552 10260
rect 17500 10217 17509 10251
rect 17509 10217 17543 10251
rect 17543 10217 17552 10251
rect 17500 10208 17552 10217
rect 7932 10072 7984 10124
rect 8392 10072 8444 10124
rect 11336 10115 11388 10124
rect 11336 10081 11345 10115
rect 11345 10081 11379 10115
rect 11379 10081 11388 10115
rect 11336 10072 11388 10081
rect 2044 10047 2096 10056
rect 2044 10013 2053 10047
rect 2053 10013 2087 10047
rect 2087 10013 2096 10047
rect 2044 10004 2096 10013
rect 4160 10004 4212 10056
rect 7196 10004 7248 10056
rect 7656 10004 7708 10056
rect 10324 10047 10376 10056
rect 10324 10013 10333 10047
rect 10333 10013 10367 10047
rect 10367 10013 10376 10047
rect 10324 10004 10376 10013
rect 10876 10004 10928 10056
rect 15200 10072 15252 10124
rect 16856 10115 16908 10124
rect 16856 10081 16865 10115
rect 16865 10081 16899 10115
rect 16899 10081 16908 10115
rect 16856 10072 16908 10081
rect 6368 9936 6420 9988
rect 11612 9979 11664 9988
rect 11612 9945 11621 9979
rect 11621 9945 11655 9979
rect 11655 9945 11664 9979
rect 11612 9936 11664 9945
rect 11704 9936 11756 9988
rect 13176 10004 13228 10056
rect 13360 10004 13412 10056
rect 13452 10047 13504 10056
rect 13452 10013 13461 10047
rect 13461 10013 13495 10047
rect 13495 10013 13504 10047
rect 13452 10004 13504 10013
rect 13728 10047 13780 10056
rect 13728 10013 13737 10047
rect 13737 10013 13771 10047
rect 13771 10013 13780 10047
rect 13728 10004 13780 10013
rect 14004 10004 14056 10056
rect 16672 10004 16724 10056
rect 1860 9911 1912 9920
rect 1860 9877 1869 9911
rect 1869 9877 1903 9911
rect 1903 9877 1912 9911
rect 1860 9868 1912 9877
rect 2688 9911 2740 9920
rect 2688 9877 2697 9911
rect 2697 9877 2731 9911
rect 2731 9877 2740 9911
rect 2688 9868 2740 9877
rect 7748 9911 7800 9920
rect 7748 9877 7757 9911
rect 7757 9877 7791 9911
rect 7791 9877 7800 9911
rect 7748 9868 7800 9877
rect 13820 9868 13872 9920
rect 14464 9911 14516 9920
rect 14464 9877 14473 9911
rect 14473 9877 14507 9911
rect 14507 9877 14516 9911
rect 14464 9868 14516 9877
rect 3737 9766 3789 9818
rect 3801 9766 3853 9818
rect 3865 9766 3917 9818
rect 3929 9766 3981 9818
rect 3993 9766 4045 9818
rect 7992 9766 8044 9818
rect 8056 9766 8108 9818
rect 8120 9766 8172 9818
rect 8184 9766 8236 9818
rect 8248 9766 8300 9818
rect 12247 9766 12299 9818
rect 12311 9766 12363 9818
rect 12375 9766 12427 9818
rect 12439 9766 12491 9818
rect 12503 9766 12555 9818
rect 16502 9766 16554 9818
rect 16566 9766 16618 9818
rect 16630 9766 16682 9818
rect 16694 9766 16746 9818
rect 16758 9766 16810 9818
rect 2044 9664 2096 9716
rect 7932 9664 7984 9716
rect 2964 9596 3016 9648
rect 3608 9528 3660 9580
rect 2596 9460 2648 9512
rect 2780 9503 2832 9512
rect 2780 9469 2789 9503
rect 2789 9469 2823 9503
rect 2823 9469 2832 9503
rect 2780 9460 2832 9469
rect 2872 9503 2924 9512
rect 2872 9469 2881 9503
rect 2881 9469 2915 9503
rect 2915 9469 2924 9503
rect 2872 9460 2924 9469
rect 2136 9392 2188 9444
rect 1768 9324 1820 9376
rect 4712 9392 4764 9444
rect 6368 9639 6420 9648
rect 6368 9605 6377 9639
rect 6377 9605 6411 9639
rect 6411 9605 6420 9639
rect 6368 9596 6420 9605
rect 6276 9528 6328 9580
rect 7564 9596 7616 9648
rect 6920 9460 6972 9512
rect 7012 9503 7064 9512
rect 7012 9469 7021 9503
rect 7021 9469 7055 9503
rect 7055 9469 7064 9503
rect 7012 9460 7064 9469
rect 7840 9528 7892 9580
rect 8576 9528 8628 9580
rect 8208 9503 8260 9512
rect 8208 9469 8217 9503
rect 8217 9469 8251 9503
rect 8251 9469 8260 9503
rect 8208 9460 8260 9469
rect 8484 9503 8536 9512
rect 8484 9469 8493 9503
rect 8493 9469 8527 9503
rect 8527 9469 8536 9503
rect 8484 9460 8536 9469
rect 8852 9528 8904 9580
rect 9128 9528 9180 9580
rect 9496 9596 9548 9648
rect 13268 9707 13320 9716
rect 13268 9673 13277 9707
rect 13277 9673 13311 9707
rect 13311 9673 13320 9707
rect 13268 9664 13320 9673
rect 13452 9707 13504 9716
rect 13452 9673 13461 9707
rect 13461 9673 13495 9707
rect 13495 9673 13504 9707
rect 13452 9664 13504 9673
rect 10784 9571 10836 9580
rect 10784 9537 10793 9571
rect 10793 9537 10827 9571
rect 10827 9537 10836 9571
rect 10784 9528 10836 9537
rect 11428 9528 11480 9580
rect 11980 9528 12032 9580
rect 12808 9596 12860 9648
rect 14556 9639 14608 9648
rect 14556 9605 14574 9639
rect 14574 9605 14608 9639
rect 14556 9596 14608 9605
rect 15384 9528 15436 9580
rect 6184 9392 6236 9444
rect 9036 9392 9088 9444
rect 4160 9324 4212 9376
rect 4988 9367 5040 9376
rect 4988 9333 4997 9367
rect 4997 9333 5031 9367
rect 5031 9333 5040 9367
rect 4988 9324 5040 9333
rect 6552 9324 6604 9376
rect 7196 9324 7248 9376
rect 7932 9324 7984 9376
rect 10048 9460 10100 9512
rect 11244 9460 11296 9512
rect 11888 9503 11940 9512
rect 11888 9469 11897 9503
rect 11897 9469 11931 9503
rect 11931 9469 11940 9503
rect 11888 9460 11940 9469
rect 15016 9460 15068 9512
rect 16304 9460 16356 9512
rect 16396 9460 16448 9512
rect 10232 9392 10284 9444
rect 11612 9392 11664 9444
rect 15660 9392 15712 9444
rect 10416 9324 10468 9376
rect 11060 9324 11112 9376
rect 12072 9367 12124 9376
rect 12072 9333 12081 9367
rect 12081 9333 12115 9367
rect 12115 9333 12124 9367
rect 12072 9324 12124 9333
rect 16488 9367 16540 9376
rect 16488 9333 16497 9367
rect 16497 9333 16531 9367
rect 16531 9333 16540 9367
rect 16488 9324 16540 9333
rect 3077 9222 3129 9274
rect 3141 9222 3193 9274
rect 3205 9222 3257 9274
rect 3269 9222 3321 9274
rect 3333 9222 3385 9274
rect 7332 9222 7384 9274
rect 7396 9222 7448 9274
rect 7460 9222 7512 9274
rect 7524 9222 7576 9274
rect 7588 9222 7640 9274
rect 11587 9222 11639 9274
rect 11651 9222 11703 9274
rect 11715 9222 11767 9274
rect 11779 9222 11831 9274
rect 11843 9222 11895 9274
rect 15842 9222 15894 9274
rect 15906 9222 15958 9274
rect 15970 9222 16022 9274
rect 16034 9222 16086 9274
rect 16098 9222 16150 9274
rect 2872 9120 2924 9172
rect 5172 9120 5224 9172
rect 6552 9163 6604 9172
rect 6552 9129 6561 9163
rect 6561 9129 6595 9163
rect 6595 9129 6604 9163
rect 6552 9120 6604 9129
rect 4344 9052 4396 9104
rect 4528 9027 4580 9036
rect 4528 8993 4537 9027
rect 4537 8993 4571 9027
rect 4571 8993 4580 9027
rect 4528 8984 4580 8993
rect 1768 8959 1820 8968
rect 1768 8925 1777 8959
rect 1777 8925 1811 8959
rect 1811 8925 1820 8959
rect 1768 8916 1820 8925
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 2136 8959 2188 8968
rect 2136 8925 2145 8959
rect 2145 8925 2179 8959
rect 2179 8925 2188 8959
rect 2136 8916 2188 8925
rect 4988 8984 5040 9036
rect 5264 8984 5316 9036
rect 5908 9027 5960 9036
rect 5908 8993 5917 9027
rect 5917 8993 5951 9027
rect 5951 8993 5960 9027
rect 5908 8984 5960 8993
rect 6092 8984 6144 9036
rect 4712 8959 4764 8968
rect 4712 8925 4721 8959
rect 4721 8925 4755 8959
rect 4755 8925 4764 8959
rect 4712 8916 4764 8925
rect 1676 8780 1728 8832
rect 2688 8848 2740 8900
rect 3516 8848 3568 8900
rect 4620 8848 4672 8900
rect 4068 8780 4120 8832
rect 4528 8780 4580 8832
rect 5816 8916 5868 8968
rect 7012 9120 7064 9172
rect 7288 9120 7340 9172
rect 8208 9120 8260 9172
rect 9128 9120 9180 9172
rect 10048 9120 10100 9172
rect 10784 9163 10836 9172
rect 10784 9129 10793 9163
rect 10793 9129 10827 9163
rect 10827 9129 10836 9163
rect 10784 9120 10836 9129
rect 11428 9163 11480 9172
rect 11428 9129 11437 9163
rect 11437 9129 11471 9163
rect 11471 9129 11480 9163
rect 11428 9120 11480 9129
rect 12624 9120 12676 9172
rect 13360 9120 13412 9172
rect 10232 9052 10284 9104
rect 12992 8984 13044 9036
rect 14556 9120 14608 9172
rect 16396 9163 16448 9172
rect 16396 9129 16405 9163
rect 16405 9129 16439 9163
rect 16439 9129 16448 9163
rect 16396 9120 16448 9129
rect 7748 8959 7800 8968
rect 7748 8925 7766 8959
rect 7766 8925 7800 8959
rect 7748 8916 7800 8925
rect 7932 8916 7984 8968
rect 9496 8959 9548 8968
rect 9496 8925 9505 8959
rect 9505 8925 9539 8959
rect 9539 8925 9548 8959
rect 9496 8916 9548 8925
rect 10048 8959 10100 8968
rect 10048 8925 10057 8959
rect 10057 8925 10091 8959
rect 10091 8925 10100 8959
rect 10048 8916 10100 8925
rect 10232 8916 10284 8968
rect 8484 8848 8536 8900
rect 8852 8848 8904 8900
rect 7656 8780 7708 8832
rect 9404 8848 9456 8900
rect 12072 8848 12124 8900
rect 14372 8916 14424 8968
rect 12624 8848 12676 8900
rect 13636 8848 13688 8900
rect 14740 8959 14792 8968
rect 14740 8925 14749 8959
rect 14749 8925 14783 8959
rect 14783 8925 14792 8959
rect 14740 8916 14792 8925
rect 9680 8780 9732 8832
rect 10508 8780 10560 8832
rect 10876 8780 10928 8832
rect 11152 8823 11204 8832
rect 11152 8789 11161 8823
rect 11161 8789 11195 8823
rect 11195 8789 11204 8823
rect 11152 8780 11204 8789
rect 11888 8780 11940 8832
rect 13176 8823 13228 8832
rect 13176 8789 13185 8823
rect 13185 8789 13219 8823
rect 13219 8789 13228 8823
rect 13176 8780 13228 8789
rect 13544 8780 13596 8832
rect 14832 8848 14884 8900
rect 15016 8959 15068 8968
rect 15016 8925 15025 8959
rect 15025 8925 15059 8959
rect 15059 8925 15068 8959
rect 15016 8916 15068 8925
rect 17224 8984 17276 9036
rect 16488 8916 16540 8968
rect 15384 8848 15436 8900
rect 15752 8848 15804 8900
rect 15568 8780 15620 8832
rect 17500 8823 17552 8832
rect 17500 8789 17509 8823
rect 17509 8789 17543 8823
rect 17543 8789 17552 8823
rect 17500 8780 17552 8789
rect 3737 8678 3789 8730
rect 3801 8678 3853 8730
rect 3865 8678 3917 8730
rect 3929 8678 3981 8730
rect 3993 8678 4045 8730
rect 7992 8678 8044 8730
rect 8056 8678 8108 8730
rect 8120 8678 8172 8730
rect 8184 8678 8236 8730
rect 8248 8678 8300 8730
rect 12247 8678 12299 8730
rect 12311 8678 12363 8730
rect 12375 8678 12427 8730
rect 12439 8678 12491 8730
rect 12503 8678 12555 8730
rect 16502 8678 16554 8730
rect 16566 8678 16618 8730
rect 16630 8678 16682 8730
rect 16694 8678 16746 8730
rect 16758 8678 16810 8730
rect 1860 8576 1912 8628
rect 3516 8576 3568 8628
rect 3608 8576 3660 8628
rect 2136 8508 2188 8560
rect 2596 8508 2648 8560
rect 5356 8576 5408 8628
rect 5816 8576 5868 8628
rect 6184 8619 6236 8628
rect 6184 8585 6193 8619
rect 6193 8585 6227 8619
rect 6227 8585 6236 8619
rect 6184 8576 6236 8585
rect 7196 8576 7248 8628
rect 7748 8576 7800 8628
rect 8392 8619 8444 8628
rect 8392 8585 8401 8619
rect 8401 8585 8435 8619
rect 8435 8585 8444 8619
rect 8392 8576 8444 8585
rect 7656 8508 7708 8560
rect 1676 8483 1728 8492
rect 1676 8449 1710 8483
rect 1710 8449 1728 8483
rect 1676 8440 1728 8449
rect 3792 8440 3844 8492
rect 4068 8440 4120 8492
rect 4712 8440 4764 8492
rect 5356 8483 5408 8492
rect 5356 8449 5390 8483
rect 5390 8449 5408 8483
rect 5356 8440 5408 8449
rect 7104 8440 7156 8492
rect 3608 8415 3660 8424
rect 3608 8381 3617 8415
rect 3617 8381 3651 8415
rect 3651 8381 3660 8415
rect 3608 8372 3660 8381
rect 4528 8415 4580 8424
rect 4528 8381 4537 8415
rect 4537 8381 4571 8415
rect 4571 8381 4580 8415
rect 4528 8372 4580 8381
rect 2596 8304 2648 8356
rect 4344 8304 4396 8356
rect 5724 8372 5776 8424
rect 6828 8372 6880 8424
rect 9680 8576 9732 8628
rect 8668 8508 8720 8560
rect 9036 8508 9088 8560
rect 10232 8508 10284 8560
rect 11980 8619 12032 8628
rect 11980 8585 11989 8619
rect 11989 8585 12023 8619
rect 12023 8585 12032 8619
rect 11980 8576 12032 8585
rect 13176 8576 13228 8628
rect 8852 8440 8904 8492
rect 9404 8440 9456 8492
rect 9496 8440 9548 8492
rect 5080 8304 5132 8356
rect 7104 8304 7156 8356
rect 7564 8304 7616 8356
rect 10048 8372 10100 8424
rect 10232 8415 10284 8424
rect 10232 8381 10241 8415
rect 10241 8381 10275 8415
rect 10275 8381 10284 8415
rect 10232 8372 10284 8381
rect 11152 8372 11204 8424
rect 10784 8304 10836 8356
rect 12164 8372 12216 8424
rect 12900 8508 12952 8560
rect 14280 8576 14332 8628
rect 14740 8576 14792 8628
rect 15660 8619 15712 8628
rect 15660 8585 15669 8619
rect 15669 8585 15703 8619
rect 15703 8585 15712 8619
rect 15660 8576 15712 8585
rect 15752 8576 15804 8628
rect 17316 8576 17368 8628
rect 13452 8508 13504 8560
rect 13728 8508 13780 8560
rect 13176 8440 13228 8492
rect 13360 8440 13412 8492
rect 13820 8440 13872 8492
rect 14372 8483 14424 8492
rect 14372 8449 14381 8483
rect 14381 8449 14415 8483
rect 14415 8449 14424 8483
rect 14372 8440 14424 8449
rect 14556 8483 14608 8492
rect 14556 8449 14565 8483
rect 14565 8449 14599 8483
rect 14599 8449 14608 8483
rect 14556 8440 14608 8449
rect 15568 8483 15620 8492
rect 6460 8236 6512 8288
rect 8760 8236 8812 8288
rect 9496 8236 9548 8288
rect 13636 8304 13688 8356
rect 14740 8372 14792 8424
rect 12072 8236 12124 8288
rect 13820 8236 13872 8288
rect 13912 8279 13964 8288
rect 13912 8245 13921 8279
rect 13921 8245 13955 8279
rect 13955 8245 13964 8279
rect 13912 8236 13964 8245
rect 14372 8304 14424 8356
rect 14924 8304 14976 8356
rect 15568 8449 15577 8483
rect 15577 8449 15611 8483
rect 15611 8449 15620 8483
rect 15568 8440 15620 8449
rect 16212 8440 16264 8492
rect 15200 8372 15252 8424
rect 15476 8372 15528 8424
rect 16948 8415 17000 8424
rect 16948 8381 16957 8415
rect 16957 8381 16991 8415
rect 16991 8381 17000 8415
rect 16948 8372 17000 8381
rect 16396 8304 16448 8356
rect 3077 8134 3129 8186
rect 3141 8134 3193 8186
rect 3205 8134 3257 8186
rect 3269 8134 3321 8186
rect 3333 8134 3385 8186
rect 7332 8134 7384 8186
rect 7396 8134 7448 8186
rect 7460 8134 7512 8186
rect 7524 8134 7576 8186
rect 7588 8134 7640 8186
rect 11587 8134 11639 8186
rect 11651 8134 11703 8186
rect 11715 8134 11767 8186
rect 11779 8134 11831 8186
rect 11843 8134 11895 8186
rect 15842 8134 15894 8186
rect 15906 8134 15958 8186
rect 15970 8134 16022 8186
rect 16034 8134 16086 8186
rect 16098 8134 16150 8186
rect 3792 8075 3844 8084
rect 3792 8041 3801 8075
rect 3801 8041 3835 8075
rect 3835 8041 3844 8075
rect 3792 8032 3844 8041
rect 10600 8032 10652 8084
rect 4988 7964 5040 8016
rect 4344 7939 4396 7948
rect 4344 7905 4353 7939
rect 4353 7905 4387 7939
rect 4387 7905 4396 7939
rect 4344 7896 4396 7905
rect 5448 7871 5500 7880
rect 5448 7837 5457 7871
rect 5457 7837 5491 7871
rect 5491 7837 5500 7871
rect 5448 7828 5500 7837
rect 5908 7828 5960 7880
rect 6644 7828 6696 7880
rect 7472 7896 7524 7948
rect 7564 7939 7616 7948
rect 7564 7905 7573 7939
rect 7573 7905 7607 7939
rect 7607 7905 7616 7939
rect 7564 7896 7616 7905
rect 7748 7964 7800 8016
rect 4160 7760 4212 7812
rect 5540 7760 5592 7812
rect 7656 7828 7708 7880
rect 12716 8032 12768 8084
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 12992 8075 13044 8084
rect 12992 8041 13001 8075
rect 13001 8041 13035 8075
rect 13035 8041 13044 8075
rect 12992 8032 13044 8041
rect 16304 8032 16356 8084
rect 13452 7871 13504 7880
rect 13452 7837 13461 7871
rect 13461 7837 13495 7871
rect 13495 7837 13504 7871
rect 13452 7828 13504 7837
rect 14556 7896 14608 7948
rect 14004 7828 14056 7880
rect 14372 7871 14424 7880
rect 14372 7837 14381 7871
rect 14381 7837 14415 7871
rect 14415 7837 14424 7871
rect 14372 7828 14424 7837
rect 5264 7735 5316 7744
rect 5264 7701 5273 7735
rect 5273 7701 5307 7735
rect 5307 7701 5316 7735
rect 5264 7692 5316 7701
rect 6552 7692 6604 7744
rect 7288 7692 7340 7744
rect 10324 7692 10376 7744
rect 11060 7692 11112 7744
rect 12808 7760 12860 7812
rect 12716 7692 12768 7744
rect 12992 7692 13044 7744
rect 14648 7692 14700 7744
rect 15016 7692 15068 7744
rect 17500 7803 17552 7812
rect 17500 7769 17518 7803
rect 17518 7769 17552 7803
rect 17500 7760 17552 7769
rect 3737 7590 3789 7642
rect 3801 7590 3853 7642
rect 3865 7590 3917 7642
rect 3929 7590 3981 7642
rect 3993 7590 4045 7642
rect 7992 7590 8044 7642
rect 8056 7590 8108 7642
rect 8120 7590 8172 7642
rect 8184 7590 8236 7642
rect 8248 7590 8300 7642
rect 12247 7590 12299 7642
rect 12311 7590 12363 7642
rect 12375 7590 12427 7642
rect 12439 7590 12491 7642
rect 12503 7590 12555 7642
rect 16502 7590 16554 7642
rect 16566 7590 16618 7642
rect 16630 7590 16682 7642
rect 16694 7590 16746 7642
rect 16758 7590 16810 7642
rect 7288 7531 7340 7540
rect 7288 7497 7297 7531
rect 7297 7497 7331 7531
rect 7331 7497 7340 7531
rect 7288 7488 7340 7497
rect 7472 7488 7524 7540
rect 10324 7488 10376 7540
rect 12716 7488 12768 7540
rect 13544 7488 13596 7540
rect 4988 7420 5040 7472
rect 7380 7463 7432 7472
rect 7380 7429 7389 7463
rect 7389 7429 7423 7463
rect 7423 7429 7432 7463
rect 7380 7420 7432 7429
rect 9588 7420 9640 7472
rect 4160 7352 4212 7404
rect 9128 7352 9180 7404
rect 9772 7352 9824 7404
rect 12072 7420 12124 7472
rect 12992 7420 13044 7472
rect 2964 7284 3016 7336
rect 4252 7327 4304 7336
rect 4252 7293 4261 7327
rect 4261 7293 4295 7327
rect 4295 7293 4304 7327
rect 4252 7284 4304 7293
rect 7656 7284 7708 7336
rect 2872 7191 2924 7200
rect 2872 7157 2881 7191
rect 2881 7157 2915 7191
rect 2915 7157 2924 7191
rect 2872 7148 2924 7157
rect 8208 7148 8260 7200
rect 11980 7395 12032 7404
rect 11980 7361 11989 7395
rect 11989 7361 12023 7395
rect 12023 7361 12032 7395
rect 11980 7352 12032 7361
rect 12164 7395 12216 7404
rect 12164 7361 12173 7395
rect 12173 7361 12207 7395
rect 12207 7361 12216 7395
rect 12164 7352 12216 7361
rect 12348 7395 12400 7404
rect 12348 7361 12357 7395
rect 12357 7361 12391 7395
rect 12391 7361 12400 7395
rect 12348 7352 12400 7361
rect 12532 7395 12584 7404
rect 12532 7361 12539 7395
rect 12539 7361 12584 7395
rect 12532 7352 12584 7361
rect 12716 7395 12768 7404
rect 12716 7361 12725 7395
rect 12725 7361 12759 7395
rect 12759 7361 12768 7395
rect 12716 7352 12768 7361
rect 12808 7395 12860 7404
rect 12808 7361 12822 7395
rect 12822 7361 12856 7395
rect 12856 7361 12860 7395
rect 12808 7352 12860 7361
rect 13084 7395 13136 7404
rect 13084 7361 13093 7395
rect 13093 7361 13127 7395
rect 13127 7361 13136 7395
rect 13084 7352 13136 7361
rect 13268 7395 13320 7404
rect 13268 7361 13275 7395
rect 13275 7361 13320 7395
rect 13268 7352 13320 7361
rect 12992 7284 13044 7336
rect 13636 7352 13688 7404
rect 14464 7488 14516 7540
rect 16304 7488 16356 7540
rect 13912 7420 13964 7472
rect 14004 7352 14056 7404
rect 15108 7352 15160 7404
rect 16396 7352 16448 7404
rect 17776 7395 17828 7404
rect 17776 7361 17785 7395
rect 17785 7361 17819 7395
rect 17819 7361 17828 7395
rect 17776 7352 17828 7361
rect 14280 7327 14332 7336
rect 14280 7293 14289 7327
rect 14289 7293 14323 7327
rect 14323 7293 14332 7327
rect 14280 7284 14332 7293
rect 14556 7284 14608 7336
rect 14648 7327 14700 7336
rect 14648 7293 14657 7327
rect 14657 7293 14691 7327
rect 14691 7293 14700 7327
rect 14648 7284 14700 7293
rect 12164 7216 12216 7268
rect 15016 7216 15068 7268
rect 10600 7191 10652 7200
rect 10600 7157 10609 7191
rect 10609 7157 10643 7191
rect 10643 7157 10652 7191
rect 10600 7148 10652 7157
rect 11152 7148 11204 7200
rect 12532 7148 12584 7200
rect 12900 7148 12952 7200
rect 13636 7148 13688 7200
rect 14188 7148 14240 7200
rect 14740 7148 14792 7200
rect 3077 7046 3129 7098
rect 3141 7046 3193 7098
rect 3205 7046 3257 7098
rect 3269 7046 3321 7098
rect 3333 7046 3385 7098
rect 7332 7046 7384 7098
rect 7396 7046 7448 7098
rect 7460 7046 7512 7098
rect 7524 7046 7576 7098
rect 7588 7046 7640 7098
rect 11587 7046 11639 7098
rect 11651 7046 11703 7098
rect 11715 7046 11767 7098
rect 11779 7046 11831 7098
rect 11843 7046 11895 7098
rect 15842 7046 15894 7098
rect 15906 7046 15958 7098
rect 15970 7046 16022 7098
rect 16034 7046 16086 7098
rect 16098 7046 16150 7098
rect 6184 6944 6236 6996
rect 7656 6944 7708 6996
rect 6000 6876 6052 6928
rect 10600 6944 10652 6996
rect 10508 6876 10560 6928
rect 12348 6944 12400 6996
rect 12992 6944 13044 6996
rect 14832 6944 14884 6996
rect 14740 6876 14792 6928
rect 4160 6783 4212 6792
rect 4160 6749 4169 6783
rect 4169 6749 4203 6783
rect 4203 6749 4212 6783
rect 4160 6740 4212 6749
rect 5264 6740 5316 6792
rect 6092 6783 6144 6792
rect 6092 6749 6099 6783
rect 6099 6749 6144 6783
rect 6092 6740 6144 6749
rect 7656 6808 7708 6860
rect 9036 6808 9088 6860
rect 2504 6672 2556 6724
rect 4528 6672 4580 6724
rect 6736 6672 6788 6724
rect 7656 6672 7708 6724
rect 4252 6604 4304 6656
rect 6828 6604 6880 6656
rect 7564 6604 7616 6656
rect 8208 6740 8260 6792
rect 9588 6740 9640 6792
rect 9956 6783 10008 6792
rect 9956 6749 9965 6783
rect 9965 6749 9999 6783
rect 9999 6749 10008 6783
rect 9956 6740 10008 6749
rect 10508 6783 10560 6792
rect 10508 6749 10517 6783
rect 10517 6749 10551 6783
rect 10551 6749 10560 6783
rect 10508 6740 10560 6749
rect 12164 6808 12216 6860
rect 14096 6808 14148 6860
rect 7840 6672 7892 6724
rect 8392 6672 8444 6724
rect 8944 6604 8996 6656
rect 9588 6647 9640 6656
rect 9588 6613 9597 6647
rect 9597 6613 9631 6647
rect 9631 6613 9640 6647
rect 9588 6604 9640 6613
rect 9772 6604 9824 6656
rect 10784 6715 10836 6724
rect 10784 6681 10793 6715
rect 10793 6681 10827 6715
rect 10827 6681 10836 6715
rect 10784 6672 10836 6681
rect 11888 6783 11940 6792
rect 11888 6749 11897 6783
rect 11897 6749 11931 6783
rect 11931 6749 11940 6783
rect 11888 6740 11940 6749
rect 14372 6740 14424 6792
rect 14464 6783 14516 6792
rect 14464 6749 14473 6783
rect 14473 6749 14507 6783
rect 14507 6749 14516 6783
rect 14464 6740 14516 6749
rect 15476 6851 15528 6860
rect 15476 6817 15485 6851
rect 15485 6817 15519 6851
rect 15519 6817 15528 6851
rect 15476 6808 15528 6817
rect 13452 6672 13504 6724
rect 14280 6672 14332 6724
rect 10968 6604 11020 6656
rect 12624 6647 12676 6656
rect 12624 6613 12633 6647
rect 12633 6613 12667 6647
rect 12667 6613 12676 6647
rect 12624 6604 12676 6613
rect 13728 6604 13780 6656
rect 15660 6647 15712 6656
rect 15660 6613 15669 6647
rect 15669 6613 15703 6647
rect 15703 6613 15712 6647
rect 15660 6604 15712 6613
rect 15752 6647 15804 6656
rect 15752 6613 15761 6647
rect 15761 6613 15795 6647
rect 15795 6613 15804 6647
rect 15752 6604 15804 6613
rect 16212 6604 16264 6656
rect 16396 6672 16448 6724
rect 16856 6672 16908 6724
rect 17500 6604 17552 6656
rect 3737 6502 3789 6554
rect 3801 6502 3853 6554
rect 3865 6502 3917 6554
rect 3929 6502 3981 6554
rect 3993 6502 4045 6554
rect 7992 6502 8044 6554
rect 8056 6502 8108 6554
rect 8120 6502 8172 6554
rect 8184 6502 8236 6554
rect 8248 6502 8300 6554
rect 12247 6502 12299 6554
rect 12311 6502 12363 6554
rect 12375 6502 12427 6554
rect 12439 6502 12491 6554
rect 12503 6502 12555 6554
rect 16502 6502 16554 6554
rect 16566 6502 16618 6554
rect 16630 6502 16682 6554
rect 16694 6502 16746 6554
rect 16758 6502 16810 6554
rect 2504 6443 2556 6452
rect 2504 6409 2513 6443
rect 2513 6409 2547 6443
rect 2547 6409 2556 6443
rect 2504 6400 2556 6409
rect 4252 6400 4304 6452
rect 4528 6443 4580 6452
rect 4528 6409 4537 6443
rect 4537 6409 4571 6443
rect 4571 6409 4580 6443
rect 4528 6400 4580 6409
rect 4988 6443 5040 6452
rect 4988 6409 4997 6443
rect 4997 6409 5031 6443
rect 5031 6409 5040 6443
rect 4988 6400 5040 6409
rect 5448 6443 5500 6452
rect 5448 6409 5457 6443
rect 5457 6409 5491 6443
rect 5491 6409 5500 6443
rect 5448 6400 5500 6409
rect 6920 6400 6972 6452
rect 7932 6400 7984 6452
rect 8254 6400 8306 6452
rect 8392 6400 8444 6452
rect 9128 6443 9180 6452
rect 9128 6409 9137 6443
rect 9137 6409 9171 6443
rect 9171 6409 9180 6443
rect 9128 6400 9180 6409
rect 10784 6400 10836 6452
rect 15660 6443 15712 6452
rect 15660 6409 15669 6443
rect 15669 6409 15703 6443
rect 15703 6409 15712 6443
rect 15660 6400 15712 6409
rect 2872 6264 2924 6316
rect 3424 6264 3476 6316
rect 4896 6264 4948 6316
rect 6552 6307 6604 6316
rect 6552 6273 6556 6307
rect 6556 6273 6590 6307
rect 6590 6273 6604 6307
rect 6552 6264 6604 6273
rect 6644 6307 6696 6316
rect 6644 6273 6653 6307
rect 6653 6273 6687 6307
rect 6687 6273 6696 6307
rect 6644 6264 6696 6273
rect 6920 6307 6972 6316
rect 6920 6273 6934 6307
rect 6934 6273 6972 6307
rect 6920 6264 6972 6273
rect 7564 6307 7616 6316
rect 7564 6273 7573 6307
rect 7573 6273 7607 6307
rect 7607 6273 7616 6307
rect 7564 6264 7616 6273
rect 7748 6264 7800 6316
rect 8944 6307 8996 6316
rect 8944 6273 8953 6307
rect 8953 6273 8987 6307
rect 8987 6273 8996 6307
rect 8944 6264 8996 6273
rect 4804 6239 4856 6248
rect 4804 6205 4813 6239
rect 4813 6205 4847 6239
rect 4847 6205 4856 6239
rect 4804 6196 4856 6205
rect 6184 6239 6236 6248
rect 6184 6205 6193 6239
rect 6193 6205 6227 6239
rect 6227 6205 6236 6239
rect 6184 6196 6236 6205
rect 7840 6196 7892 6248
rect 7932 6196 7984 6248
rect 6736 6128 6788 6180
rect 7380 6128 7432 6180
rect 9772 6128 9824 6180
rect 11060 6375 11112 6384
rect 11060 6341 11069 6375
rect 11069 6341 11103 6375
rect 11103 6341 11112 6375
rect 11060 6332 11112 6341
rect 13268 6332 13320 6384
rect 15292 6332 15344 6384
rect 15568 6332 15620 6384
rect 11152 6307 11204 6316
rect 11152 6273 11166 6307
rect 11166 6273 11200 6307
rect 11200 6273 11204 6307
rect 11152 6264 11204 6273
rect 12440 6264 12492 6316
rect 12624 6307 12676 6316
rect 12624 6273 12633 6307
rect 12633 6273 12667 6307
rect 12667 6273 12676 6307
rect 12624 6264 12676 6273
rect 15016 6307 15068 6316
rect 15016 6273 15025 6307
rect 15025 6273 15059 6307
rect 15059 6273 15068 6307
rect 15016 6264 15068 6273
rect 16304 6264 16356 6316
rect 16856 6400 16908 6452
rect 17776 6307 17828 6316
rect 17776 6273 17785 6307
rect 17785 6273 17819 6307
rect 17819 6273 17828 6307
rect 17776 6264 17828 6273
rect 11336 6196 11388 6248
rect 12256 6239 12308 6248
rect 12256 6205 12265 6239
rect 12265 6205 12299 6239
rect 12299 6205 12308 6239
rect 12256 6196 12308 6205
rect 14096 6196 14148 6248
rect 15476 6196 15528 6248
rect 15844 6239 15896 6248
rect 15844 6205 15853 6239
rect 15853 6205 15887 6239
rect 15887 6205 15896 6239
rect 15844 6196 15896 6205
rect 16396 6196 16448 6248
rect 13084 6128 13136 6180
rect 4068 6060 4120 6112
rect 6276 6060 6328 6112
rect 7288 6103 7340 6112
rect 7288 6069 7297 6103
rect 7297 6069 7331 6103
rect 7331 6069 7340 6103
rect 7288 6060 7340 6069
rect 8116 6060 8168 6112
rect 11428 6060 11480 6112
rect 3077 5958 3129 6010
rect 3141 5958 3193 6010
rect 3205 5958 3257 6010
rect 3269 5958 3321 6010
rect 3333 5958 3385 6010
rect 7332 5958 7384 6010
rect 7396 5958 7448 6010
rect 7460 5958 7512 6010
rect 7524 5958 7576 6010
rect 7588 5958 7640 6010
rect 11587 5958 11639 6010
rect 11651 5958 11703 6010
rect 11715 5958 11767 6010
rect 11779 5958 11831 6010
rect 11843 5958 11895 6010
rect 15842 5958 15894 6010
rect 15906 5958 15958 6010
rect 15970 5958 16022 6010
rect 16034 5958 16086 6010
rect 16098 5958 16150 6010
rect 4344 5856 4396 5908
rect 3424 5788 3476 5840
rect 4068 5788 4120 5840
rect 6644 5856 6696 5908
rect 4436 5763 4488 5772
rect 4436 5729 4445 5763
rect 4445 5729 4479 5763
rect 4479 5729 4488 5763
rect 4436 5720 4488 5729
rect 6184 5788 6236 5840
rect 7012 5788 7064 5840
rect 6920 5720 6972 5772
rect 11336 5856 11388 5908
rect 14924 5899 14976 5908
rect 14924 5865 14933 5899
rect 14933 5865 14967 5899
rect 14967 5865 14976 5899
rect 14924 5856 14976 5865
rect 9496 5763 9548 5772
rect 9496 5729 9505 5763
rect 9505 5729 9539 5763
rect 9539 5729 9548 5763
rect 9496 5720 9548 5729
rect 13452 5788 13504 5840
rect 15384 5788 15436 5840
rect 11060 5720 11112 5772
rect 11152 5720 11204 5772
rect 4528 5652 4580 5704
rect 5540 5695 5592 5704
rect 5540 5661 5549 5695
rect 5549 5661 5583 5695
rect 5583 5661 5592 5695
rect 5540 5652 5592 5661
rect 6276 5695 6328 5704
rect 6276 5661 6285 5695
rect 6285 5661 6319 5695
rect 6319 5661 6328 5695
rect 6276 5652 6328 5661
rect 6460 5695 6512 5704
rect 6460 5661 6469 5695
rect 6469 5661 6503 5695
rect 6503 5661 6512 5695
rect 6460 5652 6512 5661
rect 6828 5695 6880 5704
rect 6828 5661 6837 5695
rect 6837 5661 6871 5695
rect 6871 5661 6880 5695
rect 6828 5652 6880 5661
rect 7012 5695 7064 5704
rect 7012 5661 7021 5695
rect 7021 5661 7055 5695
rect 7055 5661 7064 5695
rect 7012 5652 7064 5661
rect 10968 5695 11020 5704
rect 10968 5661 10977 5695
rect 10977 5661 11011 5695
rect 11011 5661 11020 5695
rect 10968 5652 11020 5661
rect 11244 5695 11296 5704
rect 11244 5661 11253 5695
rect 11253 5661 11287 5695
rect 11287 5661 11296 5695
rect 11244 5652 11296 5661
rect 11428 5652 11480 5704
rect 7748 5584 7800 5636
rect 7840 5584 7892 5636
rect 12992 5720 13044 5772
rect 13268 5763 13320 5772
rect 13268 5729 13277 5763
rect 13277 5729 13311 5763
rect 13311 5729 13320 5763
rect 13268 5720 13320 5729
rect 13544 5720 13596 5772
rect 14372 5763 14424 5772
rect 14372 5729 14381 5763
rect 14381 5729 14415 5763
rect 14415 5729 14424 5763
rect 14372 5720 14424 5729
rect 12256 5695 12308 5704
rect 12256 5661 12265 5695
rect 12265 5661 12299 5695
rect 12299 5661 12308 5695
rect 12256 5652 12308 5661
rect 12440 5652 12492 5704
rect 15660 5720 15712 5772
rect 15844 5720 15896 5772
rect 14556 5695 14608 5704
rect 14556 5661 14565 5695
rect 14565 5661 14599 5695
rect 14599 5661 14608 5695
rect 14556 5652 14608 5661
rect 15384 5695 15436 5704
rect 15384 5661 15393 5695
rect 15393 5661 15427 5695
rect 15427 5661 15436 5695
rect 15384 5652 15436 5661
rect 17776 5763 17828 5772
rect 17776 5729 17785 5763
rect 17785 5729 17819 5763
rect 17819 5729 17828 5763
rect 17776 5720 17828 5729
rect 12716 5584 12768 5636
rect 13544 5584 13596 5636
rect 4988 5516 5040 5568
rect 6092 5559 6144 5568
rect 6092 5525 6101 5559
rect 6101 5525 6135 5559
rect 6135 5525 6144 5559
rect 6092 5516 6144 5525
rect 6276 5516 6328 5568
rect 8944 5559 8996 5568
rect 8944 5525 8953 5559
rect 8953 5525 8987 5559
rect 8987 5525 8996 5559
rect 8944 5516 8996 5525
rect 13360 5516 13412 5568
rect 15200 5559 15252 5568
rect 15200 5525 15209 5559
rect 15209 5525 15243 5559
rect 15243 5525 15252 5559
rect 15200 5516 15252 5525
rect 15752 5584 15804 5636
rect 17040 5516 17092 5568
rect 3737 5414 3789 5466
rect 3801 5414 3853 5466
rect 3865 5414 3917 5466
rect 3929 5414 3981 5466
rect 3993 5414 4045 5466
rect 7992 5414 8044 5466
rect 8056 5414 8108 5466
rect 8120 5414 8172 5466
rect 8184 5414 8236 5466
rect 8248 5414 8300 5466
rect 12247 5414 12299 5466
rect 12311 5414 12363 5466
rect 12375 5414 12427 5466
rect 12439 5414 12491 5466
rect 12503 5414 12555 5466
rect 16502 5414 16554 5466
rect 16566 5414 16618 5466
rect 16630 5414 16682 5466
rect 16694 5414 16746 5466
rect 16758 5414 16810 5466
rect 4068 5312 4120 5364
rect 7012 5312 7064 5364
rect 8944 5312 8996 5364
rect 9036 5312 9088 5364
rect 10416 5312 10468 5364
rect 10968 5312 11020 5364
rect 11060 5355 11112 5364
rect 11060 5321 11069 5355
rect 11069 5321 11103 5355
rect 11103 5321 11112 5355
rect 11060 5312 11112 5321
rect 13268 5312 13320 5364
rect 4344 5287 4396 5296
rect 2872 5219 2924 5228
rect 2872 5185 2906 5219
rect 2906 5185 2924 5219
rect 2872 5176 2924 5185
rect 4344 5253 4378 5287
rect 4378 5253 4396 5287
rect 4344 5244 4396 5253
rect 15200 5244 15252 5296
rect 4068 5151 4120 5160
rect 4068 5117 4077 5151
rect 4077 5117 4111 5151
rect 4111 5117 4120 5151
rect 4068 5108 4120 5117
rect 7288 5219 7340 5228
rect 7288 5185 7297 5219
rect 7297 5185 7331 5219
rect 7331 5185 7340 5219
rect 7288 5176 7340 5185
rect 7564 5219 7616 5228
rect 7564 5185 7573 5219
rect 7573 5185 7607 5219
rect 7607 5185 7616 5219
rect 7564 5176 7616 5185
rect 9588 5176 9640 5228
rect 11428 5176 11480 5228
rect 5540 5015 5592 5024
rect 5540 4981 5549 5015
rect 5549 4981 5583 5015
rect 5583 4981 5592 5015
rect 5540 4972 5592 4981
rect 6644 5108 6696 5160
rect 8852 5151 8904 5160
rect 8852 5117 8861 5151
rect 8861 5117 8895 5151
rect 8895 5117 8904 5151
rect 8852 5108 8904 5117
rect 9036 5151 9088 5160
rect 9036 5117 9045 5151
rect 9045 5117 9079 5151
rect 9079 5117 9088 5151
rect 9036 5108 9088 5117
rect 6828 5040 6880 5092
rect 7012 5083 7064 5092
rect 7012 5049 7021 5083
rect 7021 5049 7055 5083
rect 7055 5049 7064 5083
rect 7012 5040 7064 5049
rect 8024 5040 8076 5092
rect 9772 5108 9824 5160
rect 10140 5151 10192 5160
rect 10140 5117 10149 5151
rect 10149 5117 10183 5151
rect 10183 5117 10192 5151
rect 10140 5108 10192 5117
rect 10232 5151 10284 5160
rect 10232 5117 10266 5151
rect 10266 5117 10284 5151
rect 10232 5108 10284 5117
rect 10416 5151 10468 5160
rect 10416 5117 10425 5151
rect 10425 5117 10459 5151
rect 10459 5117 10468 5151
rect 13176 5176 13228 5228
rect 13728 5219 13780 5228
rect 13728 5185 13737 5219
rect 13737 5185 13771 5219
rect 13771 5185 13780 5219
rect 13728 5176 13780 5185
rect 13820 5219 13872 5228
rect 13820 5185 13854 5219
rect 13854 5185 13872 5219
rect 13820 5176 13872 5185
rect 14832 5176 14884 5228
rect 10416 5108 10468 5117
rect 12808 5151 12860 5160
rect 12808 5117 12817 5151
rect 12817 5117 12851 5151
rect 12851 5117 12860 5151
rect 12808 5108 12860 5117
rect 13084 5108 13136 5160
rect 14648 5108 14700 5160
rect 6920 4972 6972 5024
rect 8300 4972 8352 5024
rect 9680 5040 9732 5092
rect 12716 5040 12768 5092
rect 11336 4972 11388 5024
rect 13544 4972 13596 5024
rect 16212 4972 16264 5024
rect 17592 5015 17644 5024
rect 17592 4981 17601 5015
rect 17601 4981 17635 5015
rect 17635 4981 17644 5015
rect 17592 4972 17644 4981
rect 3077 4870 3129 4922
rect 3141 4870 3193 4922
rect 3205 4870 3257 4922
rect 3269 4870 3321 4922
rect 3333 4870 3385 4922
rect 7332 4870 7384 4922
rect 7396 4870 7448 4922
rect 7460 4870 7512 4922
rect 7524 4870 7576 4922
rect 7588 4870 7640 4922
rect 11587 4870 11639 4922
rect 11651 4870 11703 4922
rect 11715 4870 11767 4922
rect 11779 4870 11831 4922
rect 11843 4870 11895 4922
rect 15842 4870 15894 4922
rect 15906 4870 15958 4922
rect 15970 4870 16022 4922
rect 16034 4870 16086 4922
rect 16098 4870 16150 4922
rect 2872 4768 2924 4820
rect 4528 4811 4580 4820
rect 4528 4777 4537 4811
rect 4537 4777 4571 4811
rect 4571 4777 4580 4811
rect 4528 4768 4580 4777
rect 6460 4768 6512 4820
rect 6552 4768 6604 4820
rect 7012 4768 7064 4820
rect 4988 4675 5040 4684
rect 4988 4641 4997 4675
rect 4997 4641 5031 4675
rect 5031 4641 5040 4675
rect 4988 4632 5040 4641
rect 5172 4675 5224 4684
rect 5172 4641 5181 4675
rect 5181 4641 5215 4675
rect 5215 4641 5224 4675
rect 5172 4632 5224 4641
rect 5908 4632 5960 4684
rect 6736 4632 6788 4684
rect 7748 4768 7800 4820
rect 7656 4700 7708 4752
rect 10416 4768 10468 4820
rect 11152 4768 11204 4820
rect 13544 4811 13596 4820
rect 13544 4777 13553 4811
rect 13553 4777 13587 4811
rect 13587 4777 13596 4811
rect 13544 4768 13596 4777
rect 14832 4768 14884 4820
rect 15384 4768 15436 4820
rect 9496 4700 9548 4752
rect 7748 4632 7800 4684
rect 9772 4632 9824 4684
rect 9864 4675 9916 4684
rect 9864 4641 9873 4675
rect 9873 4641 9907 4675
rect 9907 4641 9916 4675
rect 9864 4632 9916 4641
rect 10232 4675 10284 4684
rect 10232 4641 10266 4675
rect 10266 4641 10284 4675
rect 10232 4632 10284 4641
rect 10416 4675 10468 4684
rect 10416 4641 10425 4675
rect 10425 4641 10459 4675
rect 10459 4641 10468 4675
rect 10416 4632 10468 4641
rect 3424 4564 3476 4616
rect 5540 4564 5592 4616
rect 6368 4564 6420 4616
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 8300 4607 8352 4616
rect 8300 4573 8309 4607
rect 8309 4573 8343 4607
rect 8343 4573 8352 4607
rect 8300 4564 8352 4573
rect 6920 4428 6972 4480
rect 7380 4428 7432 4480
rect 10140 4607 10192 4616
rect 10140 4573 10149 4607
rect 10149 4573 10183 4607
rect 10183 4573 10192 4607
rect 10140 4564 10192 4573
rect 9680 4428 9732 4480
rect 10416 4428 10468 4480
rect 13820 4632 13872 4684
rect 14188 4632 14240 4684
rect 12624 4564 12676 4616
rect 13452 4607 13504 4616
rect 13452 4573 13461 4607
rect 13461 4573 13495 4607
rect 13495 4573 13504 4607
rect 13452 4564 13504 4573
rect 13636 4564 13688 4616
rect 14464 4607 14516 4616
rect 14464 4573 14473 4607
rect 14473 4573 14507 4607
rect 14507 4573 14516 4607
rect 14464 4564 14516 4573
rect 14556 4607 14608 4616
rect 14556 4573 14565 4607
rect 14565 4573 14599 4607
rect 14599 4573 14608 4607
rect 14556 4564 14608 4573
rect 16212 4700 16264 4752
rect 15844 4632 15896 4684
rect 17684 4811 17736 4820
rect 17684 4777 17693 4811
rect 17693 4777 17727 4811
rect 17727 4777 17736 4811
rect 17684 4768 17736 4777
rect 11336 4496 11388 4548
rect 14004 4496 14056 4548
rect 14648 4496 14700 4548
rect 17040 4539 17092 4548
rect 17040 4505 17058 4539
rect 17058 4505 17092 4539
rect 17040 4496 17092 4505
rect 12716 4471 12768 4480
rect 12716 4437 12725 4471
rect 12725 4437 12759 4471
rect 12759 4437 12768 4471
rect 12716 4428 12768 4437
rect 13452 4428 13504 4480
rect 14372 4428 14424 4480
rect 15568 4428 15620 4480
rect 15660 4428 15712 4480
rect 3737 4326 3789 4378
rect 3801 4326 3853 4378
rect 3865 4326 3917 4378
rect 3929 4326 3981 4378
rect 3993 4326 4045 4378
rect 7992 4326 8044 4378
rect 8056 4326 8108 4378
rect 8120 4326 8172 4378
rect 8184 4326 8236 4378
rect 8248 4326 8300 4378
rect 12247 4326 12299 4378
rect 12311 4326 12363 4378
rect 12375 4326 12427 4378
rect 12439 4326 12491 4378
rect 12503 4326 12555 4378
rect 16502 4326 16554 4378
rect 16566 4326 16618 4378
rect 16630 4326 16682 4378
rect 16694 4326 16746 4378
rect 16758 4326 16810 4378
rect 7380 4224 7432 4276
rect 9864 4224 9916 4276
rect 11428 4224 11480 4276
rect 12716 4224 12768 4276
rect 13544 4224 13596 4276
rect 14556 4224 14608 4276
rect 15384 4224 15436 4276
rect 15844 4224 15896 4276
rect 15476 4156 15528 4208
rect 16396 4156 16448 4208
rect 4988 4088 5040 4140
rect 7748 4131 7800 4140
rect 7748 4097 7757 4131
rect 7757 4097 7791 4131
rect 7791 4097 7800 4131
rect 7748 4088 7800 4097
rect 9772 4088 9824 4140
rect 9956 4088 10008 4140
rect 10968 4088 11020 4140
rect 5540 4020 5592 4072
rect 6736 3952 6788 4004
rect 7196 3952 7248 4004
rect 4896 3884 4948 3936
rect 5816 3884 5868 3936
rect 8392 3884 8444 3936
rect 9680 4020 9732 4072
rect 10140 4020 10192 4072
rect 12716 4131 12768 4140
rect 12716 4097 12725 4131
rect 12725 4097 12759 4131
rect 12759 4097 12768 4131
rect 12716 4088 12768 4097
rect 12808 4131 12860 4140
rect 12808 4097 12817 4131
rect 12817 4097 12851 4131
rect 12851 4097 12860 4131
rect 12808 4088 12860 4097
rect 13728 4131 13780 4140
rect 13728 4097 13737 4131
rect 13737 4097 13771 4131
rect 13771 4097 13780 4131
rect 13728 4088 13780 4097
rect 13820 4131 13872 4140
rect 13820 4097 13854 4131
rect 13854 4097 13872 4131
rect 13820 4088 13872 4097
rect 14004 4131 14056 4140
rect 14004 4097 14013 4131
rect 14013 4097 14047 4131
rect 14047 4097 14056 4131
rect 14004 4088 14056 4097
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 15752 4088 15804 4140
rect 16304 4088 16356 4140
rect 17500 4131 17552 4140
rect 17500 4097 17509 4131
rect 17509 4097 17543 4131
rect 17543 4097 17552 4131
rect 17500 4088 17552 4097
rect 8668 3952 8720 4004
rect 11244 3952 11296 4004
rect 13084 4020 13136 4072
rect 13452 4063 13504 4072
rect 13452 4029 13461 4063
rect 13461 4029 13495 4063
rect 13495 4029 13504 4063
rect 13452 4020 13504 4029
rect 15660 4020 15712 4072
rect 12440 3952 12492 4004
rect 10140 3884 10192 3936
rect 10692 3884 10744 3936
rect 10968 3884 11020 3936
rect 11980 3884 12032 3936
rect 15292 3884 15344 3936
rect 3077 3782 3129 3834
rect 3141 3782 3193 3834
rect 3205 3782 3257 3834
rect 3269 3782 3321 3834
rect 3333 3782 3385 3834
rect 7332 3782 7384 3834
rect 7396 3782 7448 3834
rect 7460 3782 7512 3834
rect 7524 3782 7576 3834
rect 7588 3782 7640 3834
rect 11587 3782 11639 3834
rect 11651 3782 11703 3834
rect 11715 3782 11767 3834
rect 11779 3782 11831 3834
rect 11843 3782 11895 3834
rect 15842 3782 15894 3834
rect 15906 3782 15958 3834
rect 15970 3782 16022 3834
rect 16034 3782 16086 3834
rect 16098 3782 16150 3834
rect 7012 3680 7064 3732
rect 7104 3680 7156 3732
rect 4988 3587 5040 3596
rect 4988 3553 4997 3587
rect 4997 3553 5031 3587
rect 5031 3553 5040 3587
rect 4988 3544 5040 3553
rect 4896 3519 4948 3528
rect 4896 3485 4905 3519
rect 4905 3485 4939 3519
rect 4939 3485 4948 3519
rect 4896 3476 4948 3485
rect 7104 3587 7156 3596
rect 7104 3553 7113 3587
rect 7113 3553 7147 3587
rect 7147 3553 7156 3587
rect 7104 3544 7156 3553
rect 4160 3408 4212 3460
rect 5632 3451 5684 3460
rect 5632 3417 5666 3451
rect 5666 3417 5684 3451
rect 5632 3408 5684 3417
rect 7196 3476 7248 3528
rect 8668 3544 8720 3596
rect 8392 3519 8444 3528
rect 8392 3485 8401 3519
rect 8401 3485 8435 3519
rect 8435 3485 8444 3519
rect 8392 3476 8444 3485
rect 10600 3655 10652 3664
rect 10600 3621 10609 3655
rect 10609 3621 10643 3655
rect 10643 3621 10652 3655
rect 10600 3612 10652 3621
rect 8852 3408 8904 3460
rect 4252 3383 4304 3392
rect 4252 3349 4261 3383
rect 4261 3349 4295 3383
rect 4295 3349 4304 3383
rect 4252 3340 4304 3349
rect 4988 3340 5040 3392
rect 7748 3340 7800 3392
rect 8944 3383 8996 3392
rect 8944 3349 8953 3383
rect 8953 3349 8987 3383
rect 8987 3349 8996 3383
rect 8944 3340 8996 3349
rect 9312 3340 9364 3392
rect 10140 3587 10192 3596
rect 10140 3553 10149 3587
rect 10149 3553 10183 3587
rect 10183 3553 10192 3587
rect 10140 3544 10192 3553
rect 10416 3544 10468 3596
rect 12716 3612 12768 3664
rect 10968 3519 11020 3528
rect 10968 3485 10977 3519
rect 10977 3485 11011 3519
rect 11011 3485 11020 3519
rect 10968 3476 11020 3485
rect 11244 3544 11296 3596
rect 12440 3544 12492 3596
rect 13728 3587 13780 3596
rect 13728 3553 13737 3587
rect 13737 3553 13771 3587
rect 13771 3553 13780 3587
rect 13728 3544 13780 3553
rect 13544 3476 13596 3528
rect 14096 3519 14148 3528
rect 14096 3485 14105 3519
rect 14105 3485 14139 3519
rect 14139 3485 14148 3519
rect 14096 3476 14148 3485
rect 15292 3587 15344 3596
rect 15292 3553 15301 3587
rect 15301 3553 15335 3587
rect 15335 3553 15344 3587
rect 15292 3544 15344 3553
rect 13176 3408 13228 3460
rect 16028 3476 16080 3528
rect 17684 3451 17736 3460
rect 17684 3417 17693 3451
rect 17693 3417 17727 3451
rect 17727 3417 17736 3451
rect 17684 3408 17736 3417
rect 14280 3383 14332 3392
rect 14280 3349 14289 3383
rect 14289 3349 14323 3383
rect 14323 3349 14332 3383
rect 14280 3340 14332 3349
rect 14740 3383 14792 3392
rect 14740 3349 14749 3383
rect 14749 3349 14783 3383
rect 14783 3349 14792 3383
rect 14740 3340 14792 3349
rect 14924 3340 14976 3392
rect 15292 3340 15344 3392
rect 3737 3238 3789 3290
rect 3801 3238 3853 3290
rect 3865 3238 3917 3290
rect 3929 3238 3981 3290
rect 3993 3238 4045 3290
rect 7992 3238 8044 3290
rect 8056 3238 8108 3290
rect 8120 3238 8172 3290
rect 8184 3238 8236 3290
rect 8248 3238 8300 3290
rect 12247 3238 12299 3290
rect 12311 3238 12363 3290
rect 12375 3238 12427 3290
rect 12439 3238 12491 3290
rect 12503 3238 12555 3290
rect 16502 3238 16554 3290
rect 16566 3238 16618 3290
rect 16630 3238 16682 3290
rect 16694 3238 16746 3290
rect 16758 3238 16810 3290
rect 5540 3179 5592 3188
rect 5540 3145 5549 3179
rect 5549 3145 5583 3179
rect 5583 3145 5592 3179
rect 5540 3136 5592 3145
rect 5632 3179 5684 3188
rect 5632 3145 5641 3179
rect 5641 3145 5675 3179
rect 5675 3145 5684 3179
rect 5632 3136 5684 3145
rect 6828 3136 6880 3188
rect 9680 3136 9732 3188
rect 4252 3068 4304 3120
rect 8944 3068 8996 3120
rect 9956 3179 10008 3188
rect 9956 3145 9965 3179
rect 9965 3145 9999 3179
rect 9999 3145 10008 3179
rect 9956 3136 10008 3145
rect 12808 3136 12860 3188
rect 13176 3179 13228 3188
rect 13176 3145 13185 3179
rect 13185 3145 13219 3179
rect 13219 3145 13228 3179
rect 13176 3136 13228 3145
rect 16028 3179 16080 3188
rect 16028 3145 16037 3179
rect 16037 3145 16071 3179
rect 16071 3145 16080 3179
rect 16028 3136 16080 3145
rect 4160 3043 4212 3052
rect 4160 3009 4169 3043
rect 4169 3009 4203 3043
rect 4203 3009 4212 3043
rect 4160 3000 4212 3009
rect 5816 3043 5868 3052
rect 5816 3009 5825 3043
rect 5825 3009 5859 3043
rect 5859 3009 5868 3043
rect 5816 3000 5868 3009
rect 7656 3000 7708 3052
rect 7932 3000 7984 3052
rect 9036 3000 9088 3052
rect 10600 3000 10652 3052
rect 12624 3068 12676 3120
rect 11980 3043 12032 3052
rect 11980 3009 12014 3043
rect 12014 3009 12032 3043
rect 11980 3000 12032 3009
rect 14280 3043 14332 3052
rect 14740 3068 14792 3120
rect 14280 3009 14298 3043
rect 14298 3009 14332 3043
rect 14280 3000 14332 3009
rect 14648 3043 14700 3052
rect 14648 3009 14657 3043
rect 14657 3009 14691 3043
rect 14691 3009 14700 3043
rect 14648 3000 14700 3009
rect 9404 2796 9456 2848
rect 13636 2796 13688 2848
rect 3077 2694 3129 2746
rect 3141 2694 3193 2746
rect 3205 2694 3257 2746
rect 3269 2694 3321 2746
rect 3333 2694 3385 2746
rect 7332 2694 7384 2746
rect 7396 2694 7448 2746
rect 7460 2694 7512 2746
rect 7524 2694 7576 2746
rect 7588 2694 7640 2746
rect 11587 2694 11639 2746
rect 11651 2694 11703 2746
rect 11715 2694 11767 2746
rect 11779 2694 11831 2746
rect 11843 2694 11895 2746
rect 15842 2694 15894 2746
rect 15906 2694 15958 2746
rect 15970 2694 16022 2746
rect 16034 2694 16086 2746
rect 16098 2694 16150 2746
rect 7196 2592 7248 2644
rect 7656 2635 7708 2644
rect 7656 2601 7665 2635
rect 7665 2601 7699 2635
rect 7699 2601 7708 2635
rect 7656 2592 7708 2601
rect 10416 2635 10468 2644
rect 10416 2601 10425 2635
rect 10425 2601 10459 2635
rect 10459 2601 10468 2635
rect 10416 2592 10468 2601
rect 14096 2635 14148 2644
rect 14096 2601 14105 2635
rect 14105 2601 14139 2635
rect 14139 2601 14148 2635
rect 14096 2592 14148 2601
rect 4988 2524 5040 2576
rect 11612 2524 11664 2576
rect 13544 2524 13596 2576
rect 6828 2456 6880 2508
rect 7932 2456 7984 2508
rect 10876 2456 10928 2508
rect 12072 2456 12124 2508
rect 14924 2524 14976 2576
rect 14648 2499 14700 2508
rect 14648 2465 14657 2499
rect 14657 2465 14691 2499
rect 14691 2465 14700 2499
rect 14648 2456 14700 2465
rect 6092 2388 6144 2440
rect 6276 2388 6328 2440
rect 7840 2431 7892 2440
rect 7840 2397 7849 2431
rect 7849 2397 7883 2431
rect 7883 2397 7892 2431
rect 7840 2388 7892 2397
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 9312 2431 9364 2440
rect 9312 2397 9346 2431
rect 9346 2397 9364 2431
rect 4068 2363 4120 2372
rect 4068 2329 4077 2363
rect 4077 2329 4111 2363
rect 4111 2329 4120 2363
rect 4068 2320 4120 2329
rect 8392 2320 8444 2372
rect 9312 2388 9364 2397
rect 10324 2388 10376 2440
rect 9680 2320 9732 2372
rect 12716 2388 12768 2440
rect 12900 2388 12952 2440
rect 13176 2388 13228 2440
rect 12164 2320 12216 2372
rect 6460 2252 6512 2304
rect 7104 2252 7156 2304
rect 10968 2252 11020 2304
rect 3737 2150 3789 2202
rect 3801 2150 3853 2202
rect 3865 2150 3917 2202
rect 3929 2150 3981 2202
rect 3993 2150 4045 2202
rect 7992 2150 8044 2202
rect 8056 2150 8108 2202
rect 8120 2150 8172 2202
rect 8184 2150 8236 2202
rect 8248 2150 8300 2202
rect 12247 2150 12299 2202
rect 12311 2150 12363 2202
rect 12375 2150 12427 2202
rect 12439 2150 12491 2202
rect 12503 2150 12555 2202
rect 16502 2150 16554 2202
rect 16566 2150 16618 2202
rect 16630 2150 16682 2202
rect 16694 2150 16746 2202
rect 16758 2150 16810 2202
<< metal2 >>
rect 9034 20613 9090 21413
rect 9678 20613 9734 21413
rect 10322 20613 10378 21413
rect 12898 20754 12954 21413
rect 12636 20726 12954 20754
rect 3077 19068 3385 19077
rect 3077 19066 3083 19068
rect 3139 19066 3163 19068
rect 3219 19066 3243 19068
rect 3299 19066 3323 19068
rect 3379 19066 3385 19068
rect 3139 19014 3141 19066
rect 3321 19014 3323 19066
rect 3077 19012 3083 19014
rect 3139 19012 3163 19014
rect 3219 19012 3243 19014
rect 3299 19012 3323 19014
rect 3379 19012 3385 19014
rect 3077 19003 3385 19012
rect 7332 19068 7640 19077
rect 7332 19066 7338 19068
rect 7394 19066 7418 19068
rect 7474 19066 7498 19068
rect 7554 19066 7578 19068
rect 7634 19066 7640 19068
rect 7394 19014 7396 19066
rect 7576 19014 7578 19066
rect 7332 19012 7338 19014
rect 7394 19012 7418 19014
rect 7474 19012 7498 19014
rect 7554 19012 7578 19014
rect 7634 19012 7640 19014
rect 7332 19003 7640 19012
rect 9048 18766 9076 20613
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 7840 18760 7892 18766
rect 7840 18702 7892 18708
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 9036 18760 9088 18766
rect 9036 18702 9088 18708
rect 9312 18760 9364 18766
rect 9312 18702 9364 18708
rect 6736 18624 6788 18630
rect 6736 18566 6788 18572
rect 3737 18524 4045 18533
rect 3737 18522 3743 18524
rect 3799 18522 3823 18524
rect 3879 18522 3903 18524
rect 3959 18522 3983 18524
rect 4039 18522 4045 18524
rect 3799 18470 3801 18522
rect 3981 18470 3983 18522
rect 3737 18468 3743 18470
rect 3799 18468 3823 18470
rect 3879 18468 3903 18470
rect 3959 18468 3983 18470
rect 4039 18468 4045 18470
rect 3737 18459 4045 18468
rect 6748 18290 6776 18566
rect 6736 18284 6788 18290
rect 6736 18226 6788 18232
rect 3077 17980 3385 17989
rect 3077 17978 3083 17980
rect 3139 17978 3163 17980
rect 3219 17978 3243 17980
rect 3299 17978 3323 17980
rect 3379 17978 3385 17980
rect 3139 17926 3141 17978
rect 3321 17926 3323 17978
rect 3077 17924 3083 17926
rect 3139 17924 3163 17926
rect 3219 17924 3243 17926
rect 3299 17924 3323 17926
rect 3379 17924 3385 17926
rect 3077 17915 3385 17924
rect 7116 17882 7144 18702
rect 7656 18624 7708 18630
rect 7656 18566 7708 18572
rect 7748 18624 7800 18630
rect 7748 18566 7800 18572
rect 7668 18426 7696 18566
rect 7656 18420 7708 18426
rect 7656 18362 7708 18368
rect 7760 18306 7788 18566
rect 7668 18278 7788 18306
rect 7332 17980 7640 17989
rect 7332 17978 7338 17980
rect 7394 17978 7418 17980
rect 7474 17978 7498 17980
rect 7554 17978 7578 17980
rect 7634 17978 7640 17980
rect 7394 17926 7396 17978
rect 7576 17926 7578 17978
rect 7332 17924 7338 17926
rect 7394 17924 7418 17926
rect 7474 17924 7498 17926
rect 7554 17924 7578 17926
rect 7634 17924 7640 17926
rect 7332 17915 7640 17924
rect 7104 17876 7156 17882
rect 7104 17818 7156 17824
rect 5172 17740 5224 17746
rect 5172 17682 5224 17688
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 5080 17672 5132 17678
rect 5080 17614 5132 17620
rect 4436 17604 4488 17610
rect 4436 17546 4488 17552
rect 4160 17536 4212 17542
rect 4160 17478 4212 17484
rect 3737 17436 4045 17445
rect 3737 17434 3743 17436
rect 3799 17434 3823 17436
rect 3879 17434 3903 17436
rect 3959 17434 3983 17436
rect 4039 17434 4045 17436
rect 3799 17382 3801 17434
rect 3981 17382 3983 17434
rect 3737 17380 3743 17382
rect 3799 17380 3823 17382
rect 3879 17380 3903 17382
rect 3959 17380 3983 17382
rect 4039 17380 4045 17382
rect 3737 17371 4045 17380
rect 2872 17196 2924 17202
rect 2872 17138 2924 17144
rect 2884 16794 2912 17138
rect 2964 16992 3016 16998
rect 2964 16934 3016 16940
rect 2872 16788 2924 16794
rect 2872 16730 2924 16736
rect 2504 16652 2556 16658
rect 2504 16594 2556 16600
rect 846 16552 902 16561
rect 846 16487 848 16496
rect 900 16487 902 16496
rect 848 16458 900 16464
rect 2516 15570 2544 16594
rect 2976 16114 3004 16934
rect 3077 16892 3385 16901
rect 3077 16890 3083 16892
rect 3139 16890 3163 16892
rect 3219 16890 3243 16892
rect 3299 16890 3323 16892
rect 3379 16890 3385 16892
rect 3139 16838 3141 16890
rect 3321 16838 3323 16890
rect 3077 16836 3083 16838
rect 3139 16836 3163 16838
rect 3219 16836 3243 16838
rect 3299 16836 3323 16838
rect 3379 16836 3385 16838
rect 3077 16827 3385 16836
rect 4172 16590 4200 17478
rect 4448 16658 4476 17546
rect 4724 17338 4752 17614
rect 4896 17536 4948 17542
rect 4896 17478 4948 17484
rect 4712 17332 4764 17338
rect 4712 17274 4764 17280
rect 4908 17270 4936 17478
rect 4896 17264 4948 17270
rect 4896 17206 4948 17212
rect 5092 16794 5120 17614
rect 5080 16788 5132 16794
rect 5080 16730 5132 16736
rect 5184 16658 5212 17682
rect 7668 17678 7696 18278
rect 7748 18216 7800 18222
rect 7748 18158 7800 18164
rect 7760 17678 7788 18158
rect 7852 17882 7880 18702
rect 8484 18692 8536 18698
rect 8484 18634 8536 18640
rect 7992 18524 8300 18533
rect 7992 18522 7998 18524
rect 8054 18522 8078 18524
rect 8134 18522 8158 18524
rect 8214 18522 8238 18524
rect 8294 18522 8300 18524
rect 8054 18470 8056 18522
rect 8236 18470 8238 18522
rect 7992 18468 7998 18470
rect 8054 18468 8078 18470
rect 8134 18468 8158 18470
rect 8214 18468 8238 18470
rect 8294 18468 8300 18470
rect 7992 18459 8300 18468
rect 7840 17876 7892 17882
rect 7840 17818 7892 17824
rect 8392 17808 8444 17814
rect 8392 17750 8444 17756
rect 5632 17672 5684 17678
rect 5632 17614 5684 17620
rect 7656 17672 7708 17678
rect 7656 17614 7708 17620
rect 7748 17672 7800 17678
rect 7748 17614 7800 17620
rect 5264 17332 5316 17338
rect 5264 17274 5316 17280
rect 4436 16652 4488 16658
rect 4436 16594 4488 16600
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4252 16584 4304 16590
rect 4252 16526 4304 16532
rect 3737 16348 4045 16357
rect 3737 16346 3743 16348
rect 3799 16346 3823 16348
rect 3879 16346 3903 16348
rect 3959 16346 3983 16348
rect 4039 16346 4045 16348
rect 3799 16294 3801 16346
rect 3981 16294 3983 16346
rect 3737 16292 3743 16294
rect 3799 16292 3823 16294
rect 3879 16292 3903 16294
rect 3959 16292 3983 16294
rect 4039 16292 4045 16294
rect 3737 16283 4045 16292
rect 2964 16108 3016 16114
rect 2964 16050 3016 16056
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 2504 15564 2556 15570
rect 2504 15506 2556 15512
rect 1492 15360 1544 15366
rect 1492 15302 1544 15308
rect 1504 15065 1532 15302
rect 1490 15056 1546 15065
rect 1490 14991 1546 15000
rect 1768 15020 1820 15026
rect 1768 14962 1820 14968
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 848 14544 900 14550
rect 846 14512 848 14521
rect 900 14512 902 14521
rect 846 14447 902 14456
rect 1412 13326 1440 14894
rect 1780 14618 1808 14962
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 2320 14476 2372 14482
rect 2320 14418 2372 14424
rect 1952 13932 2004 13938
rect 1952 13874 2004 13880
rect 1676 13728 1728 13734
rect 1676 13670 1728 13676
rect 1688 13326 1716 13670
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1676 13320 1728 13326
rect 1676 13262 1728 13268
rect 1030 13016 1086 13025
rect 1030 12951 1086 12960
rect 1044 12918 1072 12951
rect 1032 12912 1084 12918
rect 1032 12854 1084 12860
rect 1412 12714 1440 13262
rect 1964 12986 1992 13874
rect 1952 12980 2004 12986
rect 1952 12922 2004 12928
rect 1400 12708 1452 12714
rect 1400 12650 1452 12656
rect 1306 12336 1362 12345
rect 1306 12271 1362 12280
rect 1320 12238 1348 12271
rect 1308 12232 1360 12238
rect 1308 12174 1360 12180
rect 1412 11694 1440 12650
rect 2044 12232 2096 12238
rect 2044 12174 2096 12180
rect 1768 12096 1820 12102
rect 1768 12038 1820 12044
rect 1860 12096 1912 12102
rect 1860 12038 1912 12044
rect 1780 11830 1808 12038
rect 1768 11824 1820 11830
rect 1768 11766 1820 11772
rect 1872 11762 1900 12038
rect 1860 11756 1912 11762
rect 1860 11698 1912 11704
rect 1400 11688 1452 11694
rect 1400 11630 1452 11636
rect 1412 10674 1440 11630
rect 2056 11354 2084 12174
rect 2044 11348 2096 11354
rect 2044 11290 2096 11296
rect 2332 11218 2360 14418
rect 2516 14278 2544 15506
rect 2780 14884 2832 14890
rect 2780 14826 2832 14832
rect 2792 14414 2820 14826
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2504 14272 2556 14278
rect 2504 14214 2556 14220
rect 2516 12782 2544 14214
rect 2976 14006 3004 16050
rect 3077 15804 3385 15813
rect 3077 15802 3083 15804
rect 3139 15802 3163 15804
rect 3219 15802 3243 15804
rect 3299 15802 3323 15804
rect 3379 15802 3385 15804
rect 3139 15750 3141 15802
rect 3321 15750 3323 15802
rect 3077 15748 3083 15750
rect 3139 15748 3163 15750
rect 3219 15748 3243 15750
rect 3299 15748 3323 15750
rect 3379 15748 3385 15750
rect 3077 15739 3385 15748
rect 3436 15706 3464 16050
rect 3424 15700 3476 15706
rect 3424 15642 3476 15648
rect 4264 15570 4292 16526
rect 4436 16176 4488 16182
rect 4436 16118 4488 16124
rect 4448 15570 4476 16118
rect 5276 15978 5304 17274
rect 5644 17134 5672 17614
rect 6000 17536 6052 17542
rect 6000 17478 6052 17484
rect 6012 17202 6040 17478
rect 6000 17196 6052 17202
rect 6000 17138 6052 17144
rect 7760 17134 7788 17614
rect 7992 17436 8300 17445
rect 7992 17434 7998 17436
rect 8054 17434 8078 17436
rect 8134 17434 8158 17436
rect 8214 17434 8238 17436
rect 8294 17434 8300 17436
rect 8054 17382 8056 17434
rect 8236 17382 8238 17434
rect 7992 17380 7998 17382
rect 8054 17380 8078 17382
rect 8134 17380 8158 17382
rect 8214 17380 8238 17382
rect 8294 17380 8300 17382
rect 7992 17371 8300 17380
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 5632 17128 5684 17134
rect 5632 17070 5684 17076
rect 7748 17128 7800 17134
rect 7748 17070 7800 17076
rect 5540 16992 5592 16998
rect 5540 16934 5592 16940
rect 5552 16658 5580 16934
rect 5540 16652 5592 16658
rect 5540 16594 5592 16600
rect 5448 16448 5500 16454
rect 5448 16390 5500 16396
rect 5356 16108 5408 16114
rect 5356 16050 5408 16056
rect 5264 15972 5316 15978
rect 5264 15914 5316 15920
rect 4620 15904 4672 15910
rect 4620 15846 4672 15852
rect 4712 15904 4764 15910
rect 4712 15846 4764 15852
rect 4252 15564 4304 15570
rect 4252 15506 4304 15512
rect 4436 15564 4488 15570
rect 4436 15506 4488 15512
rect 4264 15434 4292 15506
rect 4632 15502 4660 15846
rect 4724 15706 4752 15846
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4896 15496 4948 15502
rect 4896 15438 4948 15444
rect 5172 15496 5224 15502
rect 5172 15438 5224 15444
rect 4252 15428 4304 15434
rect 4252 15370 4304 15376
rect 3737 15260 4045 15269
rect 3737 15258 3743 15260
rect 3799 15258 3823 15260
rect 3879 15258 3903 15260
rect 3959 15258 3983 15260
rect 4039 15258 4045 15260
rect 3799 15206 3801 15258
rect 3981 15206 3983 15258
rect 3737 15204 3743 15206
rect 3799 15204 3823 15206
rect 3879 15204 3903 15206
rect 3959 15204 3983 15206
rect 4039 15204 4045 15206
rect 3737 15195 4045 15204
rect 4724 15026 4752 15438
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4908 14958 4936 15438
rect 4896 14952 4948 14958
rect 4896 14894 4948 14900
rect 3516 14816 3568 14822
rect 3516 14758 3568 14764
rect 3077 14716 3385 14725
rect 3077 14714 3083 14716
rect 3139 14714 3163 14716
rect 3219 14714 3243 14716
rect 3299 14714 3323 14716
rect 3379 14714 3385 14716
rect 3139 14662 3141 14714
rect 3321 14662 3323 14714
rect 3077 14660 3083 14662
rect 3139 14660 3163 14662
rect 3219 14660 3243 14662
rect 3299 14660 3323 14662
rect 3379 14660 3385 14662
rect 3077 14651 3385 14660
rect 2964 14000 3016 14006
rect 2884 13948 2964 13954
rect 2884 13942 3016 13948
rect 2884 13926 3004 13942
rect 2688 13728 2740 13734
rect 2688 13670 2740 13676
rect 2596 13252 2648 13258
rect 2596 13194 2648 13200
rect 2504 12776 2556 12782
rect 2504 12718 2556 12724
rect 2608 12764 2636 13194
rect 2700 12986 2728 13670
rect 2780 13320 2832 13326
rect 2780 13262 2832 13268
rect 2688 12980 2740 12986
rect 2688 12922 2740 12928
rect 2688 12776 2740 12782
rect 2608 12736 2688 12764
rect 2516 12306 2544 12718
rect 2504 12300 2556 12306
rect 2504 12242 2556 12248
rect 2412 12096 2464 12102
rect 2412 12038 2464 12044
rect 2320 11212 2372 11218
rect 2320 11154 2372 11160
rect 2424 11150 2452 12038
rect 1952 11144 2004 11150
rect 1952 11086 2004 11092
rect 2412 11144 2464 11150
rect 2412 11086 2464 11092
rect 1492 11076 1544 11082
rect 1492 11018 1544 11024
rect 1504 10985 1532 11018
rect 1768 11008 1820 11014
rect 1490 10976 1546 10985
rect 1768 10950 1820 10956
rect 1490 10911 1546 10920
rect 1780 10742 1808 10950
rect 1768 10736 1820 10742
rect 1768 10678 1820 10684
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1214 10296 1270 10305
rect 1964 10266 1992 11086
rect 1214 10231 1216 10240
rect 1268 10231 1270 10240
rect 1952 10260 2004 10266
rect 1216 10202 1268 10208
rect 1952 10202 2004 10208
rect 2608 10198 2636 12736
rect 2688 12718 2740 12724
rect 2688 11008 2740 11014
rect 2688 10950 2740 10956
rect 2596 10192 2648 10198
rect 2596 10134 2648 10140
rect 2044 10056 2096 10062
rect 2044 9998 2096 10004
rect 1860 9920 1912 9926
rect 1860 9862 1912 9868
rect 1872 9625 1900 9862
rect 2056 9722 2084 9998
rect 2700 9926 2728 10950
rect 2792 10606 2820 13262
rect 2884 12714 2912 13926
rect 3424 13864 3476 13870
rect 3424 13806 3476 13812
rect 2964 13796 3016 13802
rect 2964 13738 3016 13744
rect 2976 12782 3004 13738
rect 3077 13628 3385 13637
rect 3077 13626 3083 13628
rect 3139 13626 3163 13628
rect 3219 13626 3243 13628
rect 3299 13626 3323 13628
rect 3379 13626 3385 13628
rect 3139 13574 3141 13626
rect 3321 13574 3323 13626
rect 3077 13572 3083 13574
rect 3139 13572 3163 13574
rect 3219 13572 3243 13574
rect 3299 13572 3323 13574
rect 3379 13572 3385 13574
rect 3077 13563 3385 13572
rect 3056 13524 3108 13530
rect 3056 13466 3108 13472
rect 3068 13394 3096 13466
rect 3436 13394 3464 13806
rect 3056 13388 3108 13394
rect 3056 13330 3108 13336
rect 3424 13388 3476 13394
rect 3424 13330 3476 13336
rect 3436 12986 3464 13330
rect 3528 13326 3556 14758
rect 3737 14172 4045 14181
rect 3737 14170 3743 14172
rect 3799 14170 3823 14172
rect 3879 14170 3903 14172
rect 3959 14170 3983 14172
rect 4039 14170 4045 14172
rect 3799 14118 3801 14170
rect 3981 14118 3983 14170
rect 3737 14116 3743 14118
rect 3799 14116 3823 14118
rect 3879 14116 3903 14118
rect 3959 14116 3983 14118
rect 4039 14116 4045 14118
rect 3737 14107 4045 14116
rect 4068 14000 4120 14006
rect 4068 13942 4120 13948
rect 4436 14000 4488 14006
rect 4436 13942 4488 13948
rect 4080 13394 4108 13942
rect 4068 13388 4120 13394
rect 4068 13330 4120 13336
rect 3516 13320 3568 13326
rect 3516 13262 3568 13268
rect 3424 12980 3476 12986
rect 3424 12922 3476 12928
rect 3528 12918 3556 13262
rect 3737 13084 4045 13093
rect 3737 13082 3743 13084
rect 3799 13082 3823 13084
rect 3879 13082 3903 13084
rect 3959 13082 3983 13084
rect 4039 13082 4045 13084
rect 3799 13030 3801 13082
rect 3981 13030 3983 13082
rect 3737 13028 3743 13030
rect 3799 13028 3823 13030
rect 3879 13028 3903 13030
rect 3959 13028 3983 13030
rect 4039 13028 4045 13030
rect 3737 13019 4045 13028
rect 4080 12968 4108 13330
rect 3896 12940 4108 12968
rect 3516 12912 3568 12918
rect 3516 12854 3568 12860
rect 3896 12850 3924 12940
rect 3700 12844 3752 12850
rect 3700 12786 3752 12792
rect 3884 12844 3936 12850
rect 3884 12786 3936 12792
rect 4068 12844 4120 12850
rect 4068 12786 4120 12792
rect 2964 12776 3016 12782
rect 2964 12718 3016 12724
rect 2872 12708 2924 12714
rect 2872 12650 2924 12656
rect 2872 12232 2924 12238
rect 2872 12174 2924 12180
rect 2884 11558 2912 12174
rect 2872 11552 2924 11558
rect 2872 11494 2924 11500
rect 2884 11082 2912 11494
rect 2976 11218 3004 12718
rect 3077 12540 3385 12549
rect 3077 12538 3083 12540
rect 3139 12538 3163 12540
rect 3219 12538 3243 12540
rect 3299 12538 3323 12540
rect 3379 12538 3385 12540
rect 3139 12486 3141 12538
rect 3321 12486 3323 12538
rect 3077 12484 3083 12486
rect 3139 12484 3163 12486
rect 3219 12484 3243 12486
rect 3299 12484 3323 12486
rect 3379 12484 3385 12486
rect 3077 12475 3385 12484
rect 3712 12434 3740 12786
rect 4080 12442 4108 12786
rect 4448 12646 4476 13942
rect 5184 13938 5212 15438
rect 5276 15026 5304 15914
rect 5368 15026 5396 16050
rect 5460 15570 5488 16390
rect 5552 15706 5580 16594
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5644 15366 5672 17070
rect 7332 16892 7640 16901
rect 7332 16890 7338 16892
rect 7394 16890 7418 16892
rect 7474 16890 7498 16892
rect 7554 16890 7578 16892
rect 7634 16890 7640 16892
rect 7394 16838 7396 16890
rect 7576 16838 7578 16890
rect 7332 16836 7338 16838
rect 7394 16836 7418 16838
rect 7474 16836 7498 16838
rect 7554 16836 7578 16838
rect 7634 16836 7640 16838
rect 7332 16827 7640 16836
rect 7760 16590 7788 17070
rect 6920 16584 6972 16590
rect 6920 16526 6972 16532
rect 7748 16584 7800 16590
rect 7748 16526 7800 16532
rect 5816 16108 5868 16114
rect 5816 16050 5868 16056
rect 5724 15972 5776 15978
rect 5724 15914 5776 15920
rect 5736 15502 5764 15914
rect 5828 15570 5856 16050
rect 6092 15904 6144 15910
rect 6092 15846 6144 15852
rect 5816 15564 5868 15570
rect 5816 15506 5868 15512
rect 5724 15496 5776 15502
rect 5724 15438 5776 15444
rect 5632 15360 5684 15366
rect 5632 15302 5684 15308
rect 5724 15360 5776 15366
rect 5724 15302 5776 15308
rect 5736 15178 5764 15302
rect 5460 15150 5764 15178
rect 5264 15020 5316 15026
rect 5264 14962 5316 14968
rect 5356 15020 5408 15026
rect 5356 14962 5408 14968
rect 5460 14822 5488 15150
rect 5724 14952 5776 14958
rect 5724 14894 5776 14900
rect 5448 14816 5500 14822
rect 5448 14758 5500 14764
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 4436 12640 4488 12646
rect 4436 12582 4488 12588
rect 3620 12406 3740 12434
rect 4068 12436 4120 12442
rect 3620 11762 3648 12406
rect 5184 12434 5212 13874
rect 5184 12406 5304 12434
rect 4068 12378 4120 12384
rect 4804 12300 4856 12306
rect 4804 12242 4856 12248
rect 3737 11996 4045 12005
rect 3737 11994 3743 11996
rect 3799 11994 3823 11996
rect 3879 11994 3903 11996
rect 3959 11994 3983 11996
rect 4039 11994 4045 11996
rect 3799 11942 3801 11994
rect 3981 11942 3983 11994
rect 3737 11940 3743 11942
rect 3799 11940 3823 11942
rect 3879 11940 3903 11942
rect 3959 11940 3983 11942
rect 4039 11940 4045 11942
rect 3737 11931 4045 11940
rect 4816 11898 4844 12242
rect 5172 12232 5224 12238
rect 5092 12192 5172 12220
rect 4804 11892 4856 11898
rect 4804 11834 4856 11840
rect 3608 11756 3660 11762
rect 3608 11698 3660 11704
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3077 11452 3385 11461
rect 3077 11450 3083 11452
rect 3139 11450 3163 11452
rect 3219 11450 3243 11452
rect 3299 11450 3323 11452
rect 3379 11450 3385 11452
rect 3139 11398 3141 11450
rect 3321 11398 3323 11450
rect 3077 11396 3083 11398
rect 3139 11396 3163 11398
rect 3219 11396 3243 11398
rect 3299 11396 3323 11398
rect 3379 11396 3385 11398
rect 3077 11387 3385 11396
rect 3896 11354 3924 11698
rect 4620 11620 4672 11626
rect 4620 11562 4672 11568
rect 3884 11348 3936 11354
rect 3884 11290 3936 11296
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 4632 11150 4660 11562
rect 4816 11218 4844 11834
rect 4804 11212 4856 11218
rect 4804 11154 4856 11160
rect 3056 11144 3108 11150
rect 2976 11092 3056 11098
rect 2976 11086 3108 11092
rect 4620 11144 4672 11150
rect 4620 11086 4672 11092
rect 4712 11144 4764 11150
rect 4712 11086 4764 11092
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2976 11070 3096 11086
rect 2780 10600 2832 10606
rect 2780 10542 2832 10548
rect 2688 9920 2740 9926
rect 2688 9862 2740 9868
rect 2044 9716 2096 9722
rect 2044 9658 2096 9664
rect 1858 9616 1914 9625
rect 1858 9551 1914 9560
rect 2596 9512 2648 9518
rect 2596 9454 2648 9460
rect 2700 9500 2728 9862
rect 2976 9654 3004 11070
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3240 11008 3292 11014
rect 3240 10950 3292 10956
rect 3160 10810 3188 10950
rect 3252 10810 3280 10950
rect 3737 10908 4045 10917
rect 3737 10906 3743 10908
rect 3799 10906 3823 10908
rect 3879 10906 3903 10908
rect 3959 10906 3983 10908
rect 4039 10906 4045 10908
rect 3799 10854 3801 10906
rect 3981 10854 3983 10906
rect 3737 10852 3743 10854
rect 3799 10852 3823 10854
rect 3879 10852 3903 10854
rect 3959 10852 3983 10854
rect 4039 10852 4045 10854
rect 3737 10843 4045 10852
rect 3148 10804 3200 10810
rect 3148 10746 3200 10752
rect 3240 10804 3292 10810
rect 3240 10746 3292 10752
rect 3160 10674 3188 10746
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3077 10364 3385 10373
rect 3077 10362 3083 10364
rect 3139 10362 3163 10364
rect 3219 10362 3243 10364
rect 3299 10362 3323 10364
rect 3379 10362 3385 10364
rect 3139 10310 3141 10362
rect 3321 10310 3323 10362
rect 3077 10308 3083 10310
rect 3139 10308 3163 10310
rect 3219 10308 3243 10310
rect 3299 10308 3323 10310
rect 3379 10308 3385 10310
rect 3077 10299 3385 10308
rect 2964 9648 3016 9654
rect 2964 9590 3016 9596
rect 2780 9512 2832 9518
rect 2700 9472 2780 9500
rect 2136 9444 2188 9450
rect 2136 9386 2188 9392
rect 1768 9376 1820 9382
rect 1768 9318 1820 9324
rect 1780 8974 1808 9318
rect 2148 8974 2176 9386
rect 1768 8968 1820 8974
rect 1768 8910 1820 8916
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 2136 8968 2188 8974
rect 2136 8910 2188 8916
rect 1676 8832 1728 8838
rect 1676 8774 1728 8780
rect 1688 8498 1716 8774
rect 1872 8634 1900 8910
rect 1860 8628 1912 8634
rect 1860 8570 1912 8576
rect 2148 8566 2176 8910
rect 2608 8566 2636 9454
rect 2700 8906 2728 9472
rect 2780 9454 2832 9460
rect 2872 9512 2924 9518
rect 2872 9454 2924 9460
rect 2884 9178 2912 9454
rect 2872 9172 2924 9178
rect 2872 9114 2924 9120
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2136 8560 2188 8566
rect 2136 8502 2188 8508
rect 2596 8560 2648 8566
rect 2596 8502 2648 8508
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 2608 8362 2636 8502
rect 2596 8356 2648 8362
rect 2596 8298 2648 8304
rect 2976 7342 3004 9590
rect 3077 9276 3385 9285
rect 3077 9274 3083 9276
rect 3139 9274 3163 9276
rect 3219 9274 3243 9276
rect 3299 9274 3323 9276
rect 3379 9274 3385 9276
rect 3139 9222 3141 9274
rect 3321 9222 3323 9274
rect 3077 9220 3083 9222
rect 3139 9220 3163 9222
rect 3219 9220 3243 9222
rect 3299 9220 3323 9222
rect 3379 9220 3385 9222
rect 3077 9211 3385 9220
rect 3077 8188 3385 8197
rect 3077 8186 3083 8188
rect 3139 8186 3163 8188
rect 3219 8186 3243 8188
rect 3299 8186 3323 8188
rect 3379 8186 3385 8188
rect 3139 8134 3141 8186
rect 3321 8134 3323 8186
rect 3077 8132 3083 8134
rect 3139 8132 3163 8134
rect 3219 8132 3243 8134
rect 3299 8132 3323 8134
rect 3379 8132 3385 8134
rect 3077 8123 3385 8132
rect 2964 7336 3016 7342
rect 2964 7278 3016 7284
rect 2872 7200 2924 7206
rect 2872 7142 2924 7148
rect 2504 6724 2556 6730
rect 2504 6666 2556 6672
rect 2516 6458 2544 6666
rect 2504 6452 2556 6458
rect 2504 6394 2556 6400
rect 2884 6322 2912 7142
rect 3077 7100 3385 7109
rect 3077 7098 3083 7100
rect 3139 7098 3163 7100
rect 3219 7098 3243 7100
rect 3299 7098 3323 7100
rect 3379 7098 3385 7100
rect 3139 7046 3141 7098
rect 3321 7046 3323 7098
rect 3077 7044 3083 7046
rect 3139 7044 3163 7046
rect 3219 7044 3243 7046
rect 3299 7044 3323 7046
rect 3379 7044 3385 7046
rect 3077 7035 3385 7044
rect 3436 6322 3464 10542
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 4172 10062 4200 10406
rect 4160 10056 4212 10062
rect 4160 9998 4212 10004
rect 3737 9820 4045 9829
rect 3737 9818 3743 9820
rect 3799 9818 3823 9820
rect 3879 9818 3903 9820
rect 3959 9818 3983 9820
rect 4039 9818 4045 9820
rect 3799 9766 3801 9818
rect 3981 9766 3983 9818
rect 3737 9764 3743 9766
rect 3799 9764 3823 9766
rect 3879 9764 3903 9766
rect 3959 9764 3983 9766
rect 4039 9764 4045 9766
rect 3737 9755 4045 9764
rect 4724 9738 4752 11086
rect 4632 9710 4752 9738
rect 4526 9616 4582 9625
rect 3608 9580 3660 9586
rect 4526 9551 4582 9560
rect 3608 9522 3660 9528
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3528 8634 3556 8842
rect 3620 8634 3648 9522
rect 4160 9376 4212 9382
rect 4160 9318 4212 9324
rect 4068 8832 4120 8838
rect 4068 8774 4120 8780
rect 3737 8732 4045 8741
rect 3737 8730 3743 8732
rect 3799 8730 3823 8732
rect 3879 8730 3903 8732
rect 3959 8730 3983 8732
rect 4039 8730 4045 8732
rect 3799 8678 3801 8730
rect 3981 8678 3983 8730
rect 3737 8676 3743 8678
rect 3799 8676 3823 8678
rect 3879 8676 3903 8678
rect 3959 8676 3983 8678
rect 4039 8676 4045 8678
rect 3737 8667 4045 8676
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3608 8628 3660 8634
rect 3608 8570 3660 8576
rect 4080 8498 4108 8774
rect 3792 8492 3844 8498
rect 3792 8434 3844 8440
rect 4068 8492 4120 8498
rect 4068 8434 4120 8440
rect 3608 8424 3660 8430
rect 3606 8392 3608 8401
rect 3660 8392 3662 8401
rect 3606 8327 3662 8336
rect 3804 8090 3832 8434
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 4172 7818 4200 9318
rect 4344 9104 4396 9110
rect 4344 9046 4396 9052
rect 4356 8362 4384 9046
rect 4540 9042 4568 9551
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4632 8906 4660 9710
rect 4712 9444 4764 9450
rect 4712 9386 4764 9392
rect 4724 8974 4752 9386
rect 4712 8968 4764 8974
rect 4712 8910 4764 8916
rect 4620 8900 4672 8906
rect 4620 8842 4672 8848
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4540 8430 4568 8774
rect 4724 8498 4752 8910
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4528 8424 4580 8430
rect 4528 8366 4580 8372
rect 4344 8356 4396 8362
rect 4344 8298 4396 8304
rect 4356 7954 4384 8298
rect 4344 7948 4396 7954
rect 4344 7890 4396 7896
rect 4160 7812 4212 7818
rect 4160 7754 4212 7760
rect 3737 7644 4045 7653
rect 3737 7642 3743 7644
rect 3799 7642 3823 7644
rect 3879 7642 3903 7644
rect 3959 7642 3983 7644
rect 4039 7642 4045 7644
rect 3799 7590 3801 7642
rect 3981 7590 3983 7642
rect 3737 7588 3743 7590
rect 3799 7588 3823 7590
rect 3879 7588 3903 7590
rect 3959 7588 3983 7590
rect 4039 7588 4045 7590
rect 3737 7579 4045 7588
rect 4172 7410 4200 7754
rect 4160 7404 4212 7410
rect 4160 7346 4212 7352
rect 4172 6798 4200 7346
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 3737 6556 4045 6565
rect 3737 6554 3743 6556
rect 3799 6554 3823 6556
rect 3879 6554 3903 6556
rect 3959 6554 3983 6556
rect 4039 6554 4045 6556
rect 3799 6502 3801 6554
rect 3981 6502 3983 6554
rect 3737 6500 3743 6502
rect 3799 6500 3823 6502
rect 3879 6500 3903 6502
rect 3959 6500 3983 6502
rect 4039 6500 4045 6502
rect 3737 6491 4045 6500
rect 2872 6316 2924 6322
rect 2872 6258 2924 6264
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 3077 6012 3385 6021
rect 3077 6010 3083 6012
rect 3139 6010 3163 6012
rect 3219 6010 3243 6012
rect 3299 6010 3323 6012
rect 3379 6010 3385 6012
rect 3139 5958 3141 6010
rect 3321 5958 3323 6010
rect 3077 5956 3083 5958
rect 3139 5956 3163 5958
rect 3219 5956 3243 5958
rect 3299 5956 3323 5958
rect 3379 5956 3385 5958
rect 3077 5947 3385 5956
rect 4080 5846 4108 6054
rect 3424 5840 3476 5846
rect 3424 5782 3476 5788
rect 4068 5840 4120 5846
rect 4068 5782 4120 5788
rect 2872 5228 2924 5234
rect 2872 5170 2924 5176
rect 2884 4826 2912 5170
rect 3077 4924 3385 4933
rect 3077 4922 3083 4924
rect 3139 4922 3163 4924
rect 3219 4922 3243 4924
rect 3299 4922 3323 4924
rect 3379 4922 3385 4924
rect 3139 4870 3141 4922
rect 3321 4870 3323 4922
rect 3077 4868 3083 4870
rect 3139 4868 3163 4870
rect 3219 4868 3243 4870
rect 3299 4868 3323 4870
rect 3379 4868 3385 4870
rect 3077 4859 3385 4868
rect 2872 4820 2924 4826
rect 2872 4762 2924 4768
rect 3436 4622 3464 5782
rect 3737 5468 4045 5477
rect 3737 5466 3743 5468
rect 3799 5466 3823 5468
rect 3879 5466 3903 5468
rect 3959 5466 3983 5468
rect 4039 5466 4045 5468
rect 3799 5414 3801 5466
rect 3981 5414 3983 5466
rect 3737 5412 3743 5414
rect 3799 5412 3823 5414
rect 3879 5412 3903 5414
rect 3959 5412 3983 5414
rect 4039 5412 4045 5414
rect 3737 5403 4045 5412
rect 4080 5370 4108 5782
rect 4068 5364 4120 5370
rect 4068 5306 4120 5312
rect 4068 5160 4120 5166
rect 4172 5148 4200 6734
rect 4264 6662 4292 7278
rect 4434 6896 4490 6905
rect 4434 6831 4490 6840
rect 4252 6656 4304 6662
rect 4252 6598 4304 6604
rect 4264 6458 4292 6598
rect 4252 6452 4304 6458
rect 4252 6394 4304 6400
rect 4344 5908 4396 5914
rect 4344 5850 4396 5856
rect 4356 5302 4384 5850
rect 4448 5778 4476 6831
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 4540 6458 4568 6666
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4816 6254 4844 11154
rect 5092 11150 5120 12192
rect 5172 12174 5224 12180
rect 5080 11144 5132 11150
rect 5080 11086 5132 11092
rect 4988 9376 5040 9382
rect 4988 9318 5040 9324
rect 5000 9042 5028 9318
rect 4988 9036 5040 9042
rect 4988 8978 5040 8984
rect 5092 8362 5120 11086
rect 5276 10674 5304 12406
rect 5460 12238 5488 14758
rect 5540 13728 5592 13734
rect 5540 13670 5592 13676
rect 5552 12986 5580 13670
rect 5736 13462 5764 14894
rect 6104 14618 6132 15846
rect 6644 15360 6696 15366
rect 6644 15302 6696 15308
rect 6656 15026 6684 15302
rect 6552 15020 6604 15026
rect 6552 14962 6604 14968
rect 6644 15020 6696 15026
rect 6644 14962 6696 14968
rect 6184 14816 6236 14822
rect 6184 14758 6236 14764
rect 6368 14816 6420 14822
rect 6368 14758 6420 14764
rect 6196 14618 6224 14758
rect 6092 14612 6144 14618
rect 6092 14554 6144 14560
rect 6184 14612 6236 14618
rect 6184 14554 6236 14560
rect 6380 14550 6408 14758
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 6276 14408 6328 14414
rect 6276 14350 6328 14356
rect 5724 13456 5776 13462
rect 5724 13398 5776 13404
rect 5998 13424 6054 13433
rect 5540 12980 5592 12986
rect 5540 12922 5592 12928
rect 5552 12306 5580 12922
rect 5736 12850 5764 13398
rect 5998 13359 6054 13368
rect 6012 13326 6040 13359
rect 6000 13320 6052 13326
rect 6000 13262 6052 13268
rect 5816 13184 5868 13190
rect 5816 13126 5868 13132
rect 5828 12918 5856 13126
rect 6288 12986 6316 14350
rect 6564 14074 6592 14962
rect 6932 14958 6960 16526
rect 7196 16516 7248 16522
rect 7196 16458 7248 16464
rect 7208 16250 7236 16458
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7852 16046 7880 17138
rect 8404 17134 8432 17750
rect 8496 17542 8524 18634
rect 8588 18086 8616 18702
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8576 18080 8628 18086
rect 8576 18022 8628 18028
rect 8576 17740 8628 17746
rect 8576 17682 8628 17688
rect 8668 17740 8720 17746
rect 8668 17682 8720 17688
rect 8588 17542 8616 17682
rect 8484 17536 8536 17542
rect 8484 17478 8536 17484
rect 8576 17536 8628 17542
rect 8576 17478 8628 17484
rect 8496 17202 8524 17478
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8392 17128 8444 17134
rect 8392 17070 8444 17076
rect 8680 16794 8708 17682
rect 8956 17610 8984 18566
rect 9324 18426 9352 18702
rect 9692 18426 9720 20613
rect 10336 18970 10364 20613
rect 11587 19068 11895 19077
rect 11587 19066 11593 19068
rect 11649 19066 11673 19068
rect 11729 19066 11753 19068
rect 11809 19066 11833 19068
rect 11889 19066 11895 19068
rect 11649 19014 11651 19066
rect 11831 19014 11833 19066
rect 11587 19012 11593 19014
rect 11649 19012 11673 19014
rect 11729 19012 11753 19014
rect 11809 19012 11833 19014
rect 11889 19012 11895 19014
rect 11587 19003 11895 19012
rect 12636 18970 12664 20726
rect 12898 20613 12954 20726
rect 15842 19068 16150 19077
rect 15842 19066 15848 19068
rect 15904 19066 15928 19068
rect 15984 19066 16008 19068
rect 16064 19066 16088 19068
rect 16144 19066 16150 19068
rect 15904 19014 15906 19066
rect 16086 19014 16088 19066
rect 15842 19012 15848 19014
rect 15904 19012 15928 19014
rect 15984 19012 16008 19014
rect 16064 19012 16088 19014
rect 16144 19012 16150 19014
rect 15842 19003 16150 19012
rect 10324 18964 10376 18970
rect 10324 18906 10376 18912
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 10600 18760 10652 18766
rect 10600 18702 10652 18708
rect 11152 18760 11204 18766
rect 11152 18702 11204 18708
rect 12624 18760 12676 18766
rect 12624 18702 12676 18708
rect 13084 18760 13136 18766
rect 13084 18702 13136 18708
rect 13820 18760 13872 18766
rect 13820 18702 13872 18708
rect 9772 18692 9824 18698
rect 9772 18634 9824 18640
rect 9312 18420 9364 18426
rect 9312 18362 9364 18368
rect 9680 18420 9732 18426
rect 9680 18362 9732 18368
rect 8944 17604 8996 17610
rect 8944 17546 8996 17552
rect 8668 16788 8720 16794
rect 8668 16730 8720 16736
rect 8760 16584 8812 16590
rect 8760 16526 8812 16532
rect 7992 16348 8300 16357
rect 7992 16346 7998 16348
rect 8054 16346 8078 16348
rect 8134 16346 8158 16348
rect 8214 16346 8238 16348
rect 8294 16346 8300 16348
rect 8054 16294 8056 16346
rect 8236 16294 8238 16346
rect 7992 16292 7998 16294
rect 8054 16292 8078 16294
rect 8134 16292 8158 16294
rect 8214 16292 8238 16294
rect 8294 16292 8300 16294
rect 7992 16283 8300 16292
rect 8772 16182 8800 16526
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 8944 16448 8996 16454
rect 8944 16390 8996 16396
rect 8956 16250 8984 16390
rect 9232 16250 9260 16458
rect 8944 16244 8996 16250
rect 8944 16186 8996 16192
rect 9220 16244 9272 16250
rect 9220 16186 9272 16192
rect 8760 16176 8812 16182
rect 8760 16118 8812 16124
rect 7840 16040 7892 16046
rect 7840 15982 7892 15988
rect 8944 16040 8996 16046
rect 8944 15982 8996 15988
rect 7332 15804 7640 15813
rect 7332 15802 7338 15804
rect 7394 15802 7418 15804
rect 7474 15802 7498 15804
rect 7554 15802 7578 15804
rect 7634 15802 7640 15804
rect 7394 15750 7396 15802
rect 7576 15750 7578 15802
rect 7332 15748 7338 15750
rect 7394 15748 7418 15750
rect 7474 15748 7498 15750
rect 7554 15748 7578 15750
rect 7634 15748 7640 15750
rect 7332 15739 7640 15748
rect 7104 15564 7156 15570
rect 7104 15506 7156 15512
rect 6920 14952 6972 14958
rect 6920 14894 6972 14900
rect 6932 14346 6960 14894
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6552 14068 6604 14074
rect 6552 14010 6604 14016
rect 6460 13932 6512 13938
rect 6460 13874 6512 13880
rect 6828 13932 6880 13938
rect 6828 13874 6880 13880
rect 6368 13184 6420 13190
rect 6368 13126 6420 13132
rect 6276 12980 6328 12986
rect 6276 12922 6328 12928
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 6380 12850 6408 13126
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5908 12844 5960 12850
rect 5908 12786 5960 12792
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 5632 12708 5684 12714
rect 5632 12650 5684 12656
rect 5540 12300 5592 12306
rect 5540 12242 5592 12248
rect 5448 12232 5500 12238
rect 5448 12174 5500 12180
rect 5540 11824 5592 11830
rect 5540 11766 5592 11772
rect 5356 11688 5408 11694
rect 5356 11630 5408 11636
rect 5368 11558 5396 11630
rect 5356 11552 5408 11558
rect 5356 11494 5408 11500
rect 5368 11354 5396 11494
rect 5356 11348 5408 11354
rect 5356 11290 5408 11296
rect 5264 10668 5316 10674
rect 5264 10610 5316 10616
rect 5172 9172 5224 9178
rect 5172 9114 5224 9120
rect 5080 8356 5132 8362
rect 5080 8298 5132 8304
rect 4988 8016 5040 8022
rect 4988 7958 5040 7964
rect 5000 7478 5028 7958
rect 4988 7472 5040 7478
rect 4988 7414 5040 7420
rect 4894 6760 4950 6769
rect 4894 6695 4950 6704
rect 4908 6322 4936 6695
rect 5000 6458 5028 7414
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 4896 6316 4948 6322
rect 4896 6258 4948 6264
rect 4804 6248 4856 6254
rect 4804 6190 4856 6196
rect 4436 5772 4488 5778
rect 4436 5714 4488 5720
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4120 5120 4200 5148
rect 4068 5102 4120 5108
rect 3424 4616 3476 4622
rect 3424 4558 3476 4564
rect 3737 4380 4045 4389
rect 3737 4378 3743 4380
rect 3799 4378 3823 4380
rect 3879 4378 3903 4380
rect 3959 4378 3983 4380
rect 4039 4378 4045 4380
rect 3799 4326 3801 4378
rect 3981 4326 3983 4378
rect 3737 4324 3743 4326
rect 3799 4324 3823 4326
rect 3879 4324 3903 4326
rect 3959 4324 3983 4326
rect 4039 4324 4045 4326
rect 3737 4315 4045 4324
rect 3077 3836 3385 3845
rect 3077 3834 3083 3836
rect 3139 3834 3163 3836
rect 3219 3834 3243 3836
rect 3299 3834 3323 3836
rect 3379 3834 3385 3836
rect 3139 3782 3141 3834
rect 3321 3782 3323 3834
rect 3077 3780 3083 3782
rect 3139 3780 3163 3782
rect 3219 3780 3243 3782
rect 3299 3780 3323 3782
rect 3379 3780 3385 3782
rect 3077 3771 3385 3780
rect 4172 3466 4200 5120
rect 4540 4826 4568 5646
rect 5000 5574 5028 6394
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 4528 4820 4580 4826
rect 4528 4762 4580 4768
rect 5000 4690 5028 5510
rect 5184 4729 5212 9114
rect 5276 9042 5304 10610
rect 5368 10470 5396 11290
rect 5552 11286 5580 11766
rect 5540 11280 5592 11286
rect 5540 11222 5592 11228
rect 5552 11150 5580 11222
rect 5540 11144 5592 11150
rect 5540 11086 5592 11092
rect 5540 11008 5592 11014
rect 5540 10950 5592 10956
rect 5552 10810 5580 10950
rect 5540 10804 5592 10810
rect 5540 10746 5592 10752
rect 5540 10668 5592 10674
rect 5644 10656 5672 12650
rect 5736 10674 5764 12786
rect 5920 12442 5948 12786
rect 6472 12442 6500 13874
rect 6552 13320 6604 13326
rect 6552 13262 6604 13268
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 5908 12436 5960 12442
rect 5908 12378 5960 12384
rect 6460 12436 6512 12442
rect 6564 12434 6592 13262
rect 6644 13184 6696 13190
rect 6644 13126 6696 13132
rect 6656 12714 6684 13126
rect 6644 12708 6696 12714
rect 6644 12650 6696 12656
rect 6564 12406 6684 12434
rect 6460 12378 6512 12384
rect 6092 12368 6144 12374
rect 6092 12310 6144 12316
rect 5908 11620 5960 11626
rect 5908 11562 5960 11568
rect 5816 11144 5868 11150
rect 5920 11132 5948 11562
rect 6104 11286 6132 12310
rect 6552 12232 6604 12238
rect 6552 12174 6604 12180
rect 6368 11552 6420 11558
rect 6368 11494 6420 11500
rect 6092 11280 6144 11286
rect 6092 11222 6144 11228
rect 5868 11104 5948 11132
rect 5816 11086 5868 11092
rect 5592 10628 5672 10656
rect 5724 10668 5776 10674
rect 5540 10610 5592 10616
rect 5724 10610 5776 10616
rect 5356 10464 5408 10470
rect 5356 10406 5408 10412
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 5276 8378 5304 8978
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 5368 8498 5396 8570
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 5736 8430 5764 10610
rect 5920 9042 5948 11104
rect 6000 11076 6052 11082
rect 6000 11018 6052 11024
rect 6012 10538 6040 11018
rect 6000 10532 6052 10538
rect 6000 10474 6052 10480
rect 6104 10418 6132 11222
rect 6276 11008 6328 11014
rect 6276 10950 6328 10956
rect 6012 10390 6132 10418
rect 5908 9036 5960 9042
rect 5908 8978 5960 8984
rect 5816 8968 5868 8974
rect 5816 8910 5868 8916
rect 5828 8634 5856 8910
rect 5816 8628 5868 8634
rect 5816 8570 5868 8576
rect 5724 8424 5776 8430
rect 5276 8350 5396 8378
rect 5724 8366 5776 8372
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 5276 6798 5304 7686
rect 5264 6792 5316 6798
rect 5264 6734 5316 6740
rect 5368 5137 5396 8350
rect 5448 7880 5500 7886
rect 5448 7822 5500 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 5460 6458 5488 7822
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5448 6452 5500 6458
rect 5448 6394 5500 6400
rect 5552 5710 5580 7754
rect 5540 5704 5592 5710
rect 5540 5646 5592 5652
rect 5354 5128 5410 5137
rect 5354 5063 5410 5072
rect 5540 5024 5592 5030
rect 5540 4966 5592 4972
rect 5170 4720 5226 4729
rect 4988 4684 5040 4690
rect 5170 4655 5172 4664
rect 4988 4626 5040 4632
rect 5224 4655 5226 4664
rect 5172 4626 5224 4632
rect 5000 4146 5028 4626
rect 5552 4622 5580 4966
rect 5920 4690 5948 7822
rect 6012 6934 6040 10390
rect 6288 9586 6316 10950
rect 6380 10674 6408 11494
rect 6564 11354 6592 12174
rect 6656 11762 6684 12406
rect 6748 12306 6776 13262
rect 6736 12300 6788 12306
rect 6736 12242 6788 12248
rect 6748 11762 6776 12242
rect 6644 11756 6696 11762
rect 6644 11698 6696 11704
rect 6736 11756 6788 11762
rect 6736 11698 6788 11704
rect 6552 11348 6604 11354
rect 6552 11290 6604 11296
rect 6368 10668 6420 10674
rect 6368 10610 6420 10616
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6380 9654 6408 9930
rect 6368 9648 6420 9654
rect 6368 9590 6420 9596
rect 6276 9580 6328 9586
rect 6276 9522 6328 9528
rect 6184 9444 6236 9450
rect 6184 9386 6236 9392
rect 6092 9036 6144 9042
rect 6092 8978 6144 8984
rect 6000 6928 6052 6934
rect 6000 6870 6052 6876
rect 6104 6798 6132 8978
rect 6196 8634 6224 9386
rect 6552 9376 6604 9382
rect 6552 9318 6604 9324
rect 6564 9178 6592 9318
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6184 8628 6236 8634
rect 6184 8570 6236 8576
rect 6460 8288 6512 8294
rect 6460 8230 6512 8236
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6092 6792 6144 6798
rect 6092 6734 6144 6740
rect 6104 6633 6132 6734
rect 6090 6624 6146 6633
rect 6090 6559 6146 6568
rect 6196 6254 6224 6938
rect 6184 6248 6236 6254
rect 6182 6216 6184 6225
rect 6236 6216 6238 6225
rect 6182 6151 6238 6160
rect 6196 5846 6224 6151
rect 6276 6112 6328 6118
rect 6276 6054 6328 6060
rect 6184 5840 6236 5846
rect 6184 5782 6236 5788
rect 6288 5710 6316 6054
rect 6472 5794 6500 8230
rect 6656 7886 6684 11698
rect 6840 11626 6868 13874
rect 6932 12782 6960 14282
rect 7116 14006 7144 15506
rect 7656 15496 7708 15502
rect 7656 15438 7708 15444
rect 7288 15360 7340 15366
rect 7288 15302 7340 15308
rect 7300 15094 7328 15302
rect 7288 15088 7340 15094
rect 7288 15030 7340 15036
rect 7332 14716 7640 14725
rect 7332 14714 7338 14716
rect 7394 14714 7418 14716
rect 7474 14714 7498 14716
rect 7554 14714 7578 14716
rect 7634 14714 7640 14716
rect 7394 14662 7396 14714
rect 7576 14662 7578 14714
rect 7332 14660 7338 14662
rect 7394 14660 7418 14662
rect 7474 14660 7498 14662
rect 7554 14660 7578 14662
rect 7634 14660 7640 14662
rect 7332 14651 7640 14660
rect 7668 14074 7696 15438
rect 7656 14068 7708 14074
rect 7852 14056 7880 15982
rect 8956 15570 8984 15982
rect 9232 15978 9260 16186
rect 9324 16046 9352 18362
rect 9496 18080 9548 18086
rect 9496 18022 9548 18028
rect 9508 16046 9536 18022
rect 9588 16652 9640 16658
rect 9588 16594 9640 16600
rect 9600 16114 9628 16594
rect 9588 16108 9640 16114
rect 9588 16050 9640 16056
rect 9312 16040 9364 16046
rect 9312 15982 9364 15988
rect 9496 16040 9548 16046
rect 9496 15982 9548 15988
rect 9220 15972 9272 15978
rect 9220 15914 9272 15920
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 9140 15570 9168 15846
rect 9508 15706 9536 15982
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 8944 15564 8996 15570
rect 8944 15506 8996 15512
rect 9128 15564 9180 15570
rect 9600 15552 9628 16050
rect 9680 15564 9732 15570
rect 9600 15524 9680 15552
rect 9128 15506 9180 15512
rect 9680 15506 9732 15512
rect 7992 15260 8300 15269
rect 7992 15258 7998 15260
rect 8054 15258 8078 15260
rect 8134 15258 8158 15260
rect 8214 15258 8238 15260
rect 8294 15258 8300 15260
rect 8054 15206 8056 15258
rect 8236 15206 8238 15258
rect 7992 15204 7998 15206
rect 8054 15204 8078 15206
rect 8134 15204 8158 15206
rect 8214 15204 8238 15206
rect 8294 15204 8300 15206
rect 7992 15195 8300 15204
rect 9784 15162 9812 18634
rect 9864 18624 9916 18630
rect 9864 18566 9916 18572
rect 9876 17338 9904 18566
rect 10508 18420 10560 18426
rect 10508 18362 10560 18368
rect 10140 17876 10192 17882
rect 10140 17818 10192 17824
rect 9864 17332 9916 17338
rect 9864 17274 9916 17280
rect 9956 16040 10008 16046
rect 9956 15982 10008 15988
rect 9864 15700 9916 15706
rect 9864 15642 9916 15648
rect 9876 15502 9904 15642
rect 9864 15496 9916 15502
rect 9864 15438 9916 15444
rect 9772 15156 9824 15162
rect 9772 15098 9824 15104
rect 8668 15088 8720 15094
rect 8668 15030 8720 15036
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 7992 14172 8300 14181
rect 7992 14170 7998 14172
rect 8054 14170 8078 14172
rect 8134 14170 8158 14172
rect 8214 14170 8238 14172
rect 8294 14170 8300 14172
rect 8054 14118 8056 14170
rect 8236 14118 8238 14170
rect 7992 14116 7998 14118
rect 8054 14116 8078 14118
rect 8134 14116 8158 14118
rect 8214 14116 8238 14118
rect 8294 14116 8300 14118
rect 7992 14107 8300 14116
rect 8404 14074 8432 14758
rect 8392 14068 8444 14074
rect 7852 14028 7972 14056
rect 7656 14010 7708 14016
rect 7104 14000 7156 14006
rect 7104 13942 7156 13948
rect 7944 13938 7972 14028
rect 8392 14010 8444 14016
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 7932 13932 7984 13938
rect 7932 13874 7984 13880
rect 7656 13796 7708 13802
rect 7656 13738 7708 13744
rect 7332 13628 7640 13637
rect 7332 13626 7338 13628
rect 7394 13626 7418 13628
rect 7474 13626 7498 13628
rect 7554 13626 7578 13628
rect 7634 13626 7640 13628
rect 7394 13574 7396 13626
rect 7576 13574 7578 13626
rect 7332 13572 7338 13574
rect 7394 13572 7418 13574
rect 7474 13572 7498 13574
rect 7554 13572 7578 13574
rect 7634 13572 7640 13574
rect 7332 13563 7640 13572
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6920 12776 6972 12782
rect 6920 12718 6972 12724
rect 6828 11620 6880 11626
rect 6828 11562 6880 11568
rect 6932 10742 6960 12718
rect 7024 12442 7052 12786
rect 7116 12646 7144 13262
rect 7104 12640 7156 12646
rect 7104 12582 7156 12588
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 7116 12238 7144 12582
rect 7332 12540 7640 12549
rect 7332 12538 7338 12540
rect 7394 12538 7418 12540
rect 7474 12538 7498 12540
rect 7554 12538 7578 12540
rect 7634 12538 7640 12540
rect 7394 12486 7396 12538
rect 7576 12486 7578 12538
rect 7332 12484 7338 12486
rect 7394 12484 7418 12486
rect 7474 12484 7498 12486
rect 7554 12484 7578 12486
rect 7634 12484 7640 12486
rect 7332 12475 7640 12484
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7196 12164 7248 12170
rect 7196 12106 7248 12112
rect 7012 11756 7064 11762
rect 7012 11698 7064 11704
rect 7024 11150 7052 11698
rect 7208 11150 7236 12106
rect 7332 11452 7640 11461
rect 7332 11450 7338 11452
rect 7394 11450 7418 11452
rect 7474 11450 7498 11452
rect 7554 11450 7578 11452
rect 7634 11450 7640 11452
rect 7394 11398 7396 11450
rect 7576 11398 7578 11450
rect 7332 11396 7338 11398
rect 7394 11396 7418 11398
rect 7474 11396 7498 11398
rect 7554 11396 7578 11398
rect 7634 11396 7640 11398
rect 7332 11387 7640 11396
rect 7012 11144 7064 11150
rect 7012 11086 7064 11092
rect 7196 11144 7248 11150
rect 7196 11086 7248 11092
rect 7024 10810 7052 11086
rect 7104 11008 7156 11014
rect 7104 10950 7156 10956
rect 7196 11008 7248 11014
rect 7196 10950 7248 10956
rect 7012 10804 7064 10810
rect 7012 10746 7064 10752
rect 6920 10736 6972 10742
rect 6920 10678 6972 10684
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6840 10266 6868 10610
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6920 9512 6972 9518
rect 6920 9454 6972 9460
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6932 9058 6960 9454
rect 7024 9178 7052 9454
rect 7012 9172 7064 9178
rect 7012 9114 7064 9120
rect 6932 9030 7052 9058
rect 6828 8424 6880 8430
rect 6828 8366 6880 8372
rect 6840 8294 6868 8366
rect 6840 8266 6960 8294
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6564 6322 6592 7686
rect 6736 6724 6788 6730
rect 6736 6666 6788 6672
rect 6552 6316 6604 6322
rect 6552 6258 6604 6264
rect 6644 6316 6696 6322
rect 6644 6258 6696 6264
rect 6656 5914 6684 6258
rect 6748 6186 6776 6666
rect 6828 6656 6880 6662
rect 6828 6598 6880 6604
rect 6736 6180 6788 6186
rect 6736 6122 6788 6128
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6472 5766 6592 5794
rect 6276 5704 6328 5710
rect 6276 5646 6328 5652
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 6092 5568 6144 5574
rect 6092 5510 6144 5516
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 5908 4684 5960 4690
rect 5908 4626 5960 4632
rect 5540 4616 5592 4622
rect 5540 4558 5592 4564
rect 4988 4140 5040 4146
rect 4988 4082 5040 4088
rect 4896 3936 4948 3942
rect 4896 3878 4948 3884
rect 4908 3534 4936 3878
rect 5000 3602 5028 4082
rect 5540 4072 5592 4078
rect 5540 4014 5592 4020
rect 4988 3596 5040 3602
rect 4988 3538 5040 3544
rect 4896 3528 4948 3534
rect 4896 3470 4948 3476
rect 4160 3460 4212 3466
rect 4160 3402 4212 3408
rect 3737 3292 4045 3301
rect 3737 3290 3743 3292
rect 3799 3290 3823 3292
rect 3879 3290 3903 3292
rect 3959 3290 3983 3292
rect 4039 3290 4045 3292
rect 3799 3238 3801 3290
rect 3981 3238 3983 3290
rect 3737 3236 3743 3238
rect 3799 3236 3823 3238
rect 3879 3236 3903 3238
rect 3959 3236 3983 3238
rect 4039 3236 4045 3238
rect 3737 3227 4045 3236
rect 4172 3058 4200 3402
rect 5000 3398 5028 3538
rect 4252 3392 4304 3398
rect 4252 3334 4304 3340
rect 4988 3392 5040 3398
rect 4988 3334 5040 3340
rect 4264 3126 4292 3334
rect 4252 3120 4304 3126
rect 4252 3062 4304 3068
rect 4160 3052 4212 3058
rect 4160 2994 4212 3000
rect 3077 2748 3385 2757
rect 3077 2746 3083 2748
rect 3139 2746 3163 2748
rect 3219 2746 3243 2748
rect 3299 2746 3323 2748
rect 3379 2746 3385 2748
rect 3139 2694 3141 2746
rect 3321 2694 3323 2746
rect 3077 2692 3083 2694
rect 3139 2692 3163 2694
rect 3219 2692 3243 2694
rect 3299 2692 3323 2694
rect 3379 2692 3385 2694
rect 3077 2683 3385 2692
rect 5000 2582 5028 3334
rect 5552 3194 5580 4014
rect 5816 3936 5868 3942
rect 5816 3878 5868 3884
rect 5632 3460 5684 3466
rect 5632 3402 5684 3408
rect 5644 3194 5672 3402
rect 5540 3188 5592 3194
rect 5540 3130 5592 3136
rect 5632 3188 5684 3194
rect 5632 3130 5684 3136
rect 5828 3058 5856 3878
rect 5816 3052 5868 3058
rect 5816 2994 5868 3000
rect 4988 2576 5040 2582
rect 4988 2518 5040 2524
rect 6104 2446 6132 5510
rect 6288 2446 6316 5510
rect 6472 4826 6500 5646
rect 6564 4865 6592 5766
rect 6840 5710 6868 6598
rect 6932 6458 6960 8266
rect 6920 6452 6972 6458
rect 6920 6394 6972 6400
rect 6932 6322 6960 6394
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 7024 5846 7052 9030
rect 7116 8498 7144 10950
rect 7208 10062 7236 10950
rect 7332 10364 7640 10373
rect 7332 10362 7338 10364
rect 7394 10362 7418 10364
rect 7474 10362 7498 10364
rect 7554 10362 7578 10364
rect 7634 10362 7640 10364
rect 7394 10310 7396 10362
rect 7576 10310 7578 10362
rect 7332 10308 7338 10310
rect 7394 10308 7418 10310
rect 7474 10308 7498 10310
rect 7554 10308 7578 10310
rect 7634 10308 7640 10310
rect 7332 10299 7640 10308
rect 7668 10146 7696 13738
rect 7852 12442 7880 13874
rect 7992 13084 8300 13093
rect 7992 13082 7998 13084
rect 8054 13082 8078 13084
rect 8134 13082 8158 13084
rect 8214 13082 8238 13084
rect 8294 13082 8300 13084
rect 8054 13030 8056 13082
rect 8236 13030 8238 13082
rect 7992 13028 7998 13030
rect 8054 13028 8078 13030
rect 8134 13028 8158 13030
rect 8214 13028 8238 13030
rect 8294 13028 8300 13030
rect 7992 13019 8300 13028
rect 8392 12640 8444 12646
rect 8392 12582 8444 12588
rect 7840 12436 7892 12442
rect 7840 12378 7892 12384
rect 8208 12436 8260 12442
rect 8208 12378 8260 12384
rect 7840 12300 7892 12306
rect 7840 12242 7892 12248
rect 7852 11218 7880 12242
rect 8220 12220 8248 12378
rect 8404 12374 8432 12582
rect 8392 12368 8444 12374
rect 8392 12310 8444 12316
rect 8392 12232 8444 12238
rect 8220 12192 8392 12220
rect 8392 12174 8444 12180
rect 8496 12084 8524 14962
rect 8680 14482 8708 15030
rect 9312 15020 9364 15026
rect 9312 14962 9364 14968
rect 9220 14816 9272 14822
rect 9220 14758 9272 14764
rect 8668 14476 8720 14482
rect 8668 14418 8720 14424
rect 8576 13796 8628 13802
rect 8576 13738 8628 13744
rect 8588 13258 8616 13738
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8588 12288 8616 13194
rect 8680 12434 8708 14418
rect 9232 14414 9260 14758
rect 9220 14408 9272 14414
rect 9220 14350 9272 14356
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 8772 13841 8800 14282
rect 8944 14272 8996 14278
rect 8944 14214 8996 14220
rect 8956 14006 8984 14214
rect 9324 14074 9352 14962
rect 9312 14068 9364 14074
rect 9968 14056 9996 15982
rect 10152 15910 10180 17818
rect 10232 17604 10284 17610
rect 10232 17546 10284 17552
rect 10244 17338 10272 17546
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10232 16584 10284 16590
rect 10232 16526 10284 16532
rect 10244 15978 10272 16526
rect 10232 15972 10284 15978
rect 10232 15914 10284 15920
rect 10140 15904 10192 15910
rect 10140 15846 10192 15852
rect 10324 15904 10376 15910
rect 10324 15846 10376 15852
rect 10336 15026 10364 15846
rect 10520 15162 10548 18362
rect 10612 17882 10640 18702
rect 11060 18352 11112 18358
rect 11060 18294 11112 18300
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10704 17882 10732 18226
rect 10600 17876 10652 17882
rect 10600 17818 10652 17824
rect 10692 17876 10744 17882
rect 10692 17818 10744 17824
rect 10876 17264 10928 17270
rect 10876 17206 10928 17212
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10704 16250 10732 16934
rect 10888 16590 10916 17206
rect 11072 16794 11100 18294
rect 11164 17882 11192 18702
rect 11336 18624 11388 18630
rect 11336 18566 11388 18572
rect 11428 18624 11480 18630
rect 11428 18566 11480 18572
rect 11348 18222 11376 18566
rect 11336 18216 11388 18222
rect 11336 18158 11388 18164
rect 11152 17876 11204 17882
rect 11152 17818 11204 17824
rect 11440 17678 11468 18566
rect 12247 18524 12555 18533
rect 12247 18522 12253 18524
rect 12309 18522 12333 18524
rect 12389 18522 12413 18524
rect 12469 18522 12493 18524
rect 12549 18522 12555 18524
rect 12309 18470 12311 18522
rect 12491 18470 12493 18522
rect 12247 18468 12253 18470
rect 12309 18468 12333 18470
rect 12389 18468 12413 18470
rect 12469 18468 12493 18470
rect 12549 18468 12555 18470
rect 12247 18459 12555 18468
rect 11980 18420 12032 18426
rect 11980 18362 12032 18368
rect 11587 17980 11895 17989
rect 11587 17978 11593 17980
rect 11649 17978 11673 17980
rect 11729 17978 11753 17980
rect 11809 17978 11833 17980
rect 11889 17978 11895 17980
rect 11649 17926 11651 17978
rect 11831 17926 11833 17978
rect 11587 17924 11593 17926
rect 11649 17924 11673 17926
rect 11729 17924 11753 17926
rect 11809 17924 11833 17926
rect 11889 17924 11895 17926
rect 11587 17915 11895 17924
rect 11520 17740 11572 17746
rect 11520 17682 11572 17688
rect 11428 17672 11480 17678
rect 11428 17614 11480 17620
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11060 16788 11112 16794
rect 11060 16730 11112 16736
rect 10876 16584 10928 16590
rect 10876 16526 10928 16532
rect 10600 16244 10652 16250
rect 10600 16186 10652 16192
rect 10692 16244 10744 16250
rect 10692 16186 10744 16192
rect 10612 15910 10640 16186
rect 10692 15972 10744 15978
rect 10692 15914 10744 15920
rect 10600 15904 10652 15910
rect 10600 15846 10652 15852
rect 10508 15156 10560 15162
rect 10508 15098 10560 15104
rect 10232 15020 10284 15026
rect 10232 14962 10284 14968
rect 10324 15020 10376 15026
rect 10324 14962 10376 14968
rect 10508 15020 10560 15026
rect 10508 14962 10560 14968
rect 10048 14884 10100 14890
rect 10048 14826 10100 14832
rect 10060 14074 10088 14826
rect 10244 14634 10272 14962
rect 10140 14612 10192 14618
rect 10244 14606 10456 14634
rect 10140 14554 10192 14560
rect 10152 14074 10180 14554
rect 9312 14010 9364 14016
rect 9784 14028 9996 14056
rect 10048 14068 10100 14074
rect 8944 14000 8996 14006
rect 8944 13942 8996 13948
rect 8758 13832 8814 13841
rect 8758 13767 8814 13776
rect 9680 13728 9732 13734
rect 9680 13670 9732 13676
rect 8944 13184 8996 13190
rect 8944 13126 8996 13132
rect 8680 12406 8892 12434
rect 8588 12260 8800 12288
rect 8576 12096 8628 12102
rect 8496 12056 8576 12084
rect 8576 12038 8628 12044
rect 7992 11996 8300 12005
rect 7992 11994 7998 11996
rect 8054 11994 8078 11996
rect 8134 11994 8158 11996
rect 8214 11994 8238 11996
rect 8294 11994 8300 11996
rect 8054 11942 8056 11994
rect 8236 11942 8238 11994
rect 7992 11940 7998 11942
rect 8054 11940 8078 11942
rect 8134 11940 8158 11942
rect 8214 11940 8238 11942
rect 8294 11940 8300 11942
rect 7992 11931 8300 11940
rect 8484 11552 8536 11558
rect 8484 11494 8536 11500
rect 7840 11212 7892 11218
rect 7840 11154 7892 11160
rect 7852 10554 7880 11154
rect 7992 10908 8300 10917
rect 7992 10906 7998 10908
rect 8054 10906 8078 10908
rect 8134 10906 8158 10908
rect 8214 10906 8238 10908
rect 8294 10906 8300 10908
rect 8054 10854 8056 10906
rect 8236 10854 8238 10906
rect 7992 10852 7998 10854
rect 8054 10852 8078 10854
rect 8134 10852 8158 10854
rect 8214 10852 8238 10854
rect 8294 10852 8300 10854
rect 7992 10843 8300 10852
rect 8496 10742 8524 11494
rect 8484 10736 8536 10742
rect 8484 10678 8536 10684
rect 7852 10526 7972 10554
rect 7840 10464 7892 10470
rect 7840 10406 7892 10412
rect 7576 10118 7696 10146
rect 7196 10056 7248 10062
rect 7196 9998 7248 10004
rect 7576 9654 7604 10118
rect 7656 10056 7708 10062
rect 7656 9998 7708 10004
rect 7564 9648 7616 9654
rect 7564 9590 7616 9596
rect 7196 9376 7248 9382
rect 7196 9318 7248 9324
rect 7208 8634 7236 9318
rect 7332 9276 7640 9285
rect 7332 9274 7338 9276
rect 7394 9274 7418 9276
rect 7474 9274 7498 9276
rect 7554 9274 7578 9276
rect 7634 9274 7640 9276
rect 7394 9222 7396 9274
rect 7576 9222 7578 9274
rect 7332 9220 7338 9222
rect 7394 9220 7418 9222
rect 7474 9220 7498 9222
rect 7554 9220 7578 9222
rect 7634 9220 7640 9222
rect 7332 9211 7640 9220
rect 7288 9172 7340 9178
rect 7288 9114 7340 9120
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7300 8514 7328 9114
rect 7668 8922 7696 9998
rect 7748 9920 7800 9926
rect 7748 9862 7800 9868
rect 7760 8974 7788 9862
rect 7852 9586 7880 10406
rect 7944 10130 7972 10526
rect 7932 10124 7984 10130
rect 7932 10066 7984 10072
rect 8392 10124 8444 10130
rect 8392 10066 8444 10072
rect 7992 9820 8300 9829
rect 7992 9818 7998 9820
rect 8054 9818 8078 9820
rect 8134 9818 8158 9820
rect 8214 9818 8238 9820
rect 8294 9818 8300 9820
rect 8054 9766 8056 9818
rect 8236 9766 8238 9818
rect 7992 9764 7998 9766
rect 8054 9764 8078 9766
rect 8134 9764 8158 9766
rect 8214 9764 8238 9766
rect 8294 9764 8300 9766
rect 7992 9755 8300 9764
rect 7932 9716 7984 9722
rect 7932 9658 7984 9664
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 7944 9382 7972 9658
rect 8208 9512 8260 9518
rect 8208 9454 8260 9460
rect 7932 9376 7984 9382
rect 7932 9318 7984 9324
rect 8220 9178 8248 9454
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 7104 8492 7156 8498
rect 7104 8434 7156 8440
rect 7208 8486 7328 8514
rect 7576 8894 7696 8922
rect 7748 8968 7800 8974
rect 7932 8968 7984 8974
rect 7748 8910 7800 8916
rect 7852 8916 7932 8922
rect 7852 8910 7984 8916
rect 7852 8894 7972 8910
rect 7104 8356 7156 8362
rect 7104 8298 7156 8304
rect 7012 5840 7064 5846
rect 7012 5782 7064 5788
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6828 5704 6880 5710
rect 6932 5681 6960 5714
rect 7012 5704 7064 5710
rect 6828 5646 6880 5652
rect 6918 5672 6974 5681
rect 7012 5646 7064 5652
rect 6918 5607 6974 5616
rect 7024 5370 7052 5646
rect 7012 5364 7064 5370
rect 7012 5306 7064 5312
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 7010 5128 7066 5137
rect 6550 4856 6606 4865
rect 6460 4820 6512 4826
rect 6550 4791 6552 4800
rect 6460 4762 6512 4768
rect 6604 4791 6606 4800
rect 6552 4762 6604 4768
rect 6656 4706 6684 5102
rect 6828 5092 6880 5098
rect 7010 5063 7012 5072
rect 6828 5034 6880 5040
rect 7064 5063 7066 5072
rect 7012 5034 7064 5040
rect 6472 4678 6684 4706
rect 6736 4684 6788 4690
rect 6368 4616 6420 4622
rect 6472 4604 6500 4678
rect 6736 4626 6788 4632
rect 6420 4576 6500 4604
rect 6368 4558 6420 4564
rect 6748 4010 6776 4626
rect 6840 4593 6868 5034
rect 6920 5024 6972 5030
rect 6972 4972 7052 4978
rect 6920 4966 7052 4972
rect 6932 4950 7052 4966
rect 6918 4856 6974 4865
rect 7024 4826 7052 4950
rect 6918 4791 6974 4800
rect 7012 4820 7064 4826
rect 6826 4584 6882 4593
rect 6826 4519 6882 4528
rect 6736 4004 6788 4010
rect 6736 3946 6788 3952
rect 6840 3194 6868 4519
rect 6932 4486 6960 4791
rect 7012 4762 7064 4768
rect 6920 4480 6972 4486
rect 6920 4422 6972 4428
rect 7024 3738 7052 4762
rect 7116 3738 7144 8298
rect 7208 5681 7236 8486
rect 7576 8362 7604 8894
rect 7656 8832 7708 8838
rect 7656 8774 7708 8780
rect 7668 8566 7696 8774
rect 7748 8628 7800 8634
rect 7748 8570 7800 8576
rect 7656 8560 7708 8566
rect 7656 8502 7708 8508
rect 7760 8378 7788 8570
rect 7564 8356 7616 8362
rect 7564 8298 7616 8304
rect 7668 8350 7788 8378
rect 7332 8188 7640 8197
rect 7332 8186 7338 8188
rect 7394 8186 7418 8188
rect 7474 8186 7498 8188
rect 7554 8186 7578 8188
rect 7634 8186 7640 8188
rect 7394 8134 7396 8186
rect 7576 8134 7578 8186
rect 7332 8132 7338 8134
rect 7394 8132 7418 8134
rect 7474 8132 7498 8134
rect 7554 8132 7578 8134
rect 7634 8132 7640 8134
rect 7332 8123 7640 8132
rect 7668 8072 7696 8350
rect 7576 8044 7696 8072
rect 7378 7984 7434 7993
rect 7576 7954 7604 8044
rect 7748 8016 7800 8022
rect 7748 7958 7800 7964
rect 7378 7919 7434 7928
rect 7472 7948 7524 7954
rect 7288 7744 7340 7750
rect 7288 7686 7340 7692
rect 7300 7546 7328 7686
rect 7288 7540 7340 7546
rect 7288 7482 7340 7488
rect 7392 7478 7420 7919
rect 7472 7890 7524 7896
rect 7564 7948 7616 7954
rect 7564 7890 7616 7896
rect 7484 7546 7512 7890
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7472 7540 7524 7546
rect 7472 7482 7524 7488
rect 7380 7472 7432 7478
rect 7380 7414 7432 7420
rect 7668 7342 7696 7822
rect 7656 7336 7708 7342
rect 7656 7278 7708 7284
rect 7332 7100 7640 7109
rect 7332 7098 7338 7100
rect 7394 7098 7418 7100
rect 7474 7098 7498 7100
rect 7554 7098 7578 7100
rect 7634 7098 7640 7100
rect 7394 7046 7396 7098
rect 7576 7046 7578 7098
rect 7332 7044 7338 7046
rect 7394 7044 7418 7046
rect 7474 7044 7498 7046
rect 7554 7044 7578 7046
rect 7634 7044 7640 7046
rect 7332 7035 7640 7044
rect 7668 7002 7696 7278
rect 7656 6996 7708 7002
rect 7656 6938 7708 6944
rect 7668 6866 7696 6938
rect 7656 6860 7708 6866
rect 7656 6802 7708 6808
rect 7656 6724 7708 6730
rect 7656 6666 7708 6672
rect 7564 6656 7616 6662
rect 7378 6624 7434 6633
rect 7564 6598 7616 6604
rect 7378 6559 7434 6568
rect 7286 6216 7342 6225
rect 7392 6186 7420 6559
rect 7576 6322 7604 6598
rect 7564 6316 7616 6322
rect 7564 6258 7616 6264
rect 7286 6151 7342 6160
rect 7380 6180 7432 6186
rect 7300 6118 7328 6151
rect 7380 6122 7432 6128
rect 7288 6112 7340 6118
rect 7288 6054 7340 6060
rect 7332 6012 7640 6021
rect 7332 6010 7338 6012
rect 7394 6010 7418 6012
rect 7474 6010 7498 6012
rect 7554 6010 7578 6012
rect 7634 6010 7640 6012
rect 7394 5958 7396 6010
rect 7576 5958 7578 6010
rect 7332 5956 7338 5958
rect 7394 5956 7418 5958
rect 7474 5956 7498 5958
rect 7554 5956 7578 5958
rect 7634 5956 7640 5958
rect 7332 5947 7640 5956
rect 7194 5672 7250 5681
rect 7194 5607 7250 5616
rect 7668 5522 7696 6666
rect 7760 6322 7788 7958
rect 7852 6730 7880 8894
rect 7992 8732 8300 8741
rect 7992 8730 7998 8732
rect 8054 8730 8078 8732
rect 8134 8730 8158 8732
rect 8214 8730 8238 8732
rect 8294 8730 8300 8732
rect 8054 8678 8056 8730
rect 8236 8678 8238 8730
rect 7992 8676 7998 8678
rect 8054 8676 8078 8678
rect 8134 8676 8158 8678
rect 8214 8676 8238 8678
rect 8294 8676 8300 8678
rect 7992 8667 8300 8676
rect 8404 8634 8432 10066
rect 8588 9586 8616 12038
rect 8668 11892 8720 11898
rect 8668 11834 8720 11840
rect 8680 11626 8708 11834
rect 8668 11620 8720 11626
rect 8668 11562 8720 11568
rect 8576 9580 8628 9586
rect 8576 9522 8628 9528
rect 8484 9512 8536 9518
rect 8484 9454 8536 9460
rect 8496 8906 8524 9454
rect 8484 8900 8536 8906
rect 8484 8842 8536 8848
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 7992 7644 8300 7653
rect 7992 7642 7998 7644
rect 8054 7642 8078 7644
rect 8134 7642 8158 7644
rect 8214 7642 8238 7644
rect 8294 7642 8300 7644
rect 8054 7590 8056 7642
rect 8236 7590 8238 7642
rect 7992 7588 7998 7590
rect 8054 7588 8078 7590
rect 8134 7588 8158 7590
rect 8214 7588 8238 7590
rect 8294 7588 8300 7590
rect 7992 7579 8300 7588
rect 8208 7200 8260 7206
rect 8208 7142 8260 7148
rect 8220 6798 8248 7142
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 7840 6724 7892 6730
rect 7840 6666 7892 6672
rect 8392 6724 8444 6730
rect 8392 6666 8444 6672
rect 7748 6316 7800 6322
rect 7748 6258 7800 6264
rect 7852 6254 7880 6666
rect 7992 6556 8300 6565
rect 7992 6554 7998 6556
rect 8054 6554 8078 6556
rect 8134 6554 8158 6556
rect 8214 6554 8238 6556
rect 8294 6554 8300 6556
rect 8054 6502 8056 6554
rect 8236 6502 8238 6554
rect 7992 6500 7998 6502
rect 8054 6500 8078 6502
rect 8134 6500 8158 6502
rect 8214 6500 8238 6502
rect 8294 6500 8300 6502
rect 7992 6491 8300 6500
rect 8404 6458 8432 6666
rect 7932 6452 7984 6458
rect 8254 6452 8306 6458
rect 7932 6394 7984 6400
rect 8128 6412 8254 6440
rect 7944 6254 7972 6394
rect 7840 6248 7892 6254
rect 7840 6190 7892 6196
rect 7932 6248 7984 6254
rect 7932 6190 7984 6196
rect 7852 5642 7880 6190
rect 8128 6118 8156 6412
rect 8254 6394 8306 6400
rect 8392 6452 8444 6458
rect 8392 6394 8444 6400
rect 8116 6112 8168 6118
rect 8116 6054 8168 6060
rect 7748 5636 7800 5642
rect 7748 5578 7800 5584
rect 7840 5636 7892 5642
rect 7840 5578 7892 5584
rect 7576 5494 7696 5522
rect 7576 5234 7604 5494
rect 7288 5228 7340 5234
rect 7208 5188 7288 5216
rect 7208 4010 7236 5188
rect 7288 5170 7340 5176
rect 7564 5228 7616 5234
rect 7564 5170 7616 5176
rect 7576 5114 7604 5170
rect 7576 5086 7696 5114
rect 7332 4924 7640 4933
rect 7332 4922 7338 4924
rect 7394 4922 7418 4924
rect 7474 4922 7498 4924
rect 7554 4922 7578 4924
rect 7634 4922 7640 4924
rect 7394 4870 7396 4922
rect 7576 4870 7578 4922
rect 7332 4868 7338 4870
rect 7394 4868 7418 4870
rect 7474 4868 7498 4870
rect 7554 4868 7578 4870
rect 7634 4868 7640 4870
rect 7332 4859 7640 4868
rect 7668 4758 7696 5086
rect 7760 4826 7788 5578
rect 7748 4820 7800 4826
rect 7748 4762 7800 4768
rect 7656 4752 7708 4758
rect 7656 4694 7708 4700
rect 7748 4684 7800 4690
rect 7748 4626 7800 4632
rect 7288 4616 7340 4622
rect 7286 4584 7288 4593
rect 7340 4584 7342 4593
rect 7286 4519 7342 4528
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7392 4282 7420 4422
rect 7380 4276 7432 4282
rect 7380 4218 7432 4224
rect 7760 4146 7788 4626
rect 7748 4140 7800 4146
rect 7748 4082 7800 4088
rect 7196 4004 7248 4010
rect 7196 3946 7248 3952
rect 7332 3836 7640 3845
rect 7332 3834 7338 3836
rect 7394 3834 7418 3836
rect 7474 3834 7498 3836
rect 7554 3834 7578 3836
rect 7634 3834 7640 3836
rect 7394 3782 7396 3834
rect 7576 3782 7578 3834
rect 7332 3780 7338 3782
rect 7394 3780 7418 3782
rect 7474 3780 7498 3782
rect 7554 3780 7578 3782
rect 7634 3780 7640 3782
rect 7332 3771 7640 3780
rect 7012 3732 7064 3738
rect 7012 3674 7064 3680
rect 7104 3732 7156 3738
rect 7104 3674 7156 3680
rect 7116 3602 7144 3674
rect 7104 3596 7156 3602
rect 7104 3538 7156 3544
rect 7196 3528 7248 3534
rect 7196 3470 7248 3476
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6840 2514 6868 3130
rect 7208 2650 7236 3470
rect 7748 3392 7800 3398
rect 7748 3334 7800 3340
rect 7656 3052 7708 3058
rect 7656 2994 7708 3000
rect 7332 2748 7640 2757
rect 7332 2746 7338 2748
rect 7394 2746 7418 2748
rect 7474 2746 7498 2748
rect 7554 2746 7578 2748
rect 7634 2746 7640 2748
rect 7394 2694 7396 2746
rect 7576 2694 7578 2746
rect 7332 2692 7338 2694
rect 7394 2692 7418 2694
rect 7474 2692 7498 2694
rect 7554 2692 7578 2694
rect 7634 2692 7640 2694
rect 7332 2683 7640 2692
rect 7668 2650 7696 2994
rect 7760 2774 7788 3334
rect 7852 3040 7880 5578
rect 7992 5468 8300 5477
rect 7992 5466 7998 5468
rect 8054 5466 8078 5468
rect 8134 5466 8158 5468
rect 8214 5466 8238 5468
rect 8294 5466 8300 5468
rect 8054 5414 8056 5466
rect 8236 5414 8238 5466
rect 7992 5412 7998 5414
rect 8054 5412 8078 5414
rect 8134 5412 8158 5414
rect 8214 5412 8238 5414
rect 8294 5412 8300 5414
rect 7992 5403 8300 5412
rect 8022 5128 8078 5137
rect 8022 5063 8024 5072
rect 8076 5063 8078 5072
rect 8024 5034 8076 5040
rect 8300 5024 8352 5030
rect 8300 4966 8352 4972
rect 8312 4622 8340 4966
rect 8300 4616 8352 4622
rect 8300 4558 8352 4564
rect 7992 4380 8300 4389
rect 7992 4378 7998 4380
rect 8054 4378 8078 4380
rect 8134 4378 8158 4380
rect 8214 4378 8238 4380
rect 8294 4378 8300 4380
rect 8054 4326 8056 4378
rect 8236 4326 8238 4378
rect 7992 4324 7998 4326
rect 8054 4324 8078 4326
rect 8134 4324 8158 4326
rect 8214 4324 8238 4326
rect 8294 4324 8300 4326
rect 7992 4315 8300 4324
rect 8392 3936 8444 3942
rect 8392 3878 8444 3884
rect 8404 3534 8432 3878
rect 8392 3528 8444 3534
rect 8392 3470 8444 3476
rect 7992 3292 8300 3301
rect 7992 3290 7998 3292
rect 8054 3290 8078 3292
rect 8134 3290 8158 3292
rect 8214 3290 8238 3292
rect 8294 3290 8300 3292
rect 8054 3238 8056 3290
rect 8236 3238 8238 3290
rect 7992 3236 7998 3238
rect 8054 3236 8078 3238
rect 8134 3236 8158 3238
rect 8214 3236 8238 3238
rect 8294 3236 8300 3238
rect 7992 3227 8300 3236
rect 7932 3052 7984 3058
rect 7852 3012 7932 3040
rect 7932 2994 7984 3000
rect 7760 2746 7880 2774
rect 7196 2644 7248 2650
rect 7196 2586 7248 2592
rect 7656 2644 7708 2650
rect 7656 2586 7708 2592
rect 6828 2508 6880 2514
rect 6828 2450 6880 2456
rect 7852 2446 7880 2746
rect 7944 2514 7972 2994
rect 7932 2508 7984 2514
rect 7932 2450 7984 2456
rect 8496 2446 8524 8842
rect 8680 8566 8708 11562
rect 8668 8560 8720 8566
rect 8668 8502 8720 8508
rect 8772 8294 8800 12260
rect 8864 12084 8892 12406
rect 8956 12238 8984 13126
rect 9692 12918 9720 13670
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 9220 12844 9272 12850
rect 9220 12786 9272 12792
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9232 12170 9260 12786
rect 9404 12640 9456 12646
rect 9404 12582 9456 12588
rect 9680 12640 9732 12646
rect 9680 12582 9732 12588
rect 9416 12442 9444 12582
rect 9404 12436 9456 12442
rect 9404 12378 9456 12384
rect 9220 12164 9272 12170
rect 9220 12106 9272 12112
rect 9036 12096 9088 12102
rect 8864 12056 9036 12084
rect 9036 12038 9088 12044
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8864 8906 8892 9522
rect 9048 9450 9076 12038
rect 9416 11694 9444 12378
rect 9692 12374 9720 12582
rect 9680 12368 9732 12374
rect 9680 12310 9732 12316
rect 9404 11688 9456 11694
rect 9404 11630 9456 11636
rect 9416 10810 9444 11630
rect 9784 11354 9812 14028
rect 10048 14010 10100 14016
rect 10140 14068 10192 14074
rect 10192 14028 10364 14056
rect 10140 14010 10192 14016
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 9864 13864 9916 13870
rect 9864 13806 9916 13812
rect 9876 11830 9904 13806
rect 9968 12850 9996 13874
rect 10060 13258 10088 14010
rect 10140 13456 10192 13462
rect 10140 13398 10192 13404
rect 10152 13258 10180 13398
rect 10232 13388 10284 13394
rect 10232 13330 10284 13336
rect 10048 13252 10100 13258
rect 10048 13194 10100 13200
rect 10140 13252 10192 13258
rect 10140 13194 10192 13200
rect 9956 12844 10008 12850
rect 9956 12786 10008 12792
rect 10244 12646 10272 13330
rect 10336 13326 10364 14028
rect 10324 13320 10376 13326
rect 10324 13262 10376 13268
rect 10428 12986 10456 14606
rect 10520 13530 10548 14962
rect 10704 13870 10732 15914
rect 10784 15360 10836 15366
rect 10784 15302 10836 15308
rect 10796 15026 10824 15302
rect 10784 15020 10836 15026
rect 10784 14962 10836 14968
rect 10692 13864 10744 13870
rect 10692 13806 10744 13812
rect 10508 13524 10560 13530
rect 10508 13466 10560 13472
rect 10888 13410 10916 16526
rect 10968 15020 11020 15026
rect 10968 14962 11020 14968
rect 10980 14618 11008 14962
rect 11072 14958 11100 16730
rect 11164 16182 11192 17478
rect 11336 17128 11388 17134
rect 11336 17070 11388 17076
rect 11348 16794 11376 17070
rect 11532 16946 11560 17682
rect 11440 16918 11560 16946
rect 11336 16788 11388 16794
rect 11336 16730 11388 16736
rect 11152 16176 11204 16182
rect 11204 16136 11284 16164
rect 11152 16118 11204 16124
rect 11152 15020 11204 15026
rect 11152 14962 11204 14968
rect 11060 14952 11112 14958
rect 11060 14894 11112 14900
rect 10968 14612 11020 14618
rect 10968 14554 11020 14560
rect 11072 14482 11100 14894
rect 11060 14476 11112 14482
rect 11060 14418 11112 14424
rect 11164 14074 11192 14962
rect 11152 14068 11204 14074
rect 11152 14010 11204 14016
rect 11256 13954 11284 16136
rect 11336 14476 11388 14482
rect 11336 14418 11388 14424
rect 10520 13382 10916 13410
rect 10980 13926 11284 13954
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10232 12640 10284 12646
rect 10232 12582 10284 12588
rect 9864 11824 9916 11830
rect 9864 11766 9916 11772
rect 10324 11824 10376 11830
rect 10324 11766 10376 11772
rect 9772 11348 9824 11354
rect 9772 11290 9824 11296
rect 9680 11144 9732 11150
rect 9680 11086 9732 11092
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 9494 10704 9550 10713
rect 9494 10639 9496 10648
rect 9548 10639 9550 10648
rect 9496 10610 9548 10616
rect 9692 10266 9720 11086
rect 9680 10260 9732 10266
rect 9680 10202 9732 10208
rect 9784 10198 9812 11290
rect 9772 10192 9824 10198
rect 9772 10134 9824 10140
rect 10336 10062 10364 11766
rect 10324 10056 10376 10062
rect 10324 9998 10376 10004
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 9036 9444 9088 9450
rect 9036 9386 9088 9392
rect 9140 9178 9168 9522
rect 9128 9172 9180 9178
rect 9128 9114 9180 9120
rect 9508 8974 9536 9590
rect 10048 9512 10100 9518
rect 10048 9454 10100 9460
rect 10060 9178 10088 9454
rect 10232 9444 10284 9450
rect 10232 9386 10284 9392
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10060 8974 10088 9114
rect 10244 9110 10272 9386
rect 10416 9376 10468 9382
rect 10416 9318 10468 9324
rect 10232 9104 10284 9110
rect 10232 9046 10284 9052
rect 10244 8974 10272 9046
rect 9496 8968 9548 8974
rect 9496 8910 9548 8916
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 10232 8968 10284 8974
rect 10232 8910 10284 8916
rect 8852 8900 8904 8906
rect 8852 8842 8904 8848
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 8864 8498 8892 8842
rect 9036 8560 9088 8566
rect 9036 8502 9088 8508
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8760 8288 8812 8294
rect 8760 8230 8812 8236
rect 9048 6866 9076 8502
rect 9416 8498 9444 8842
rect 9508 8498 9536 8910
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9692 8634 9720 8774
rect 9680 8628 9732 8634
rect 9680 8570 9732 8576
rect 9404 8492 9456 8498
rect 9404 8434 9456 8440
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9128 7404 9180 7410
rect 9128 7346 9180 7352
rect 9036 6860 9088 6866
rect 9036 6802 9088 6808
rect 8944 6656 8996 6662
rect 8944 6598 8996 6604
rect 8956 6322 8984 6598
rect 9140 6458 9168 7346
rect 9128 6452 9180 6458
rect 9128 6394 9180 6400
rect 8944 6316 8996 6322
rect 8944 6258 8996 6264
rect 8944 5568 8996 5574
rect 8944 5510 8996 5516
rect 8956 5370 8984 5510
rect 8944 5364 8996 5370
rect 8944 5306 8996 5312
rect 9036 5364 9088 5370
rect 9036 5306 9088 5312
rect 9048 5166 9076 5306
rect 8852 5160 8904 5166
rect 8852 5102 8904 5108
rect 9036 5160 9088 5166
rect 9036 5102 9088 5108
rect 8668 4004 8720 4010
rect 8668 3946 8720 3952
rect 8680 3602 8708 3946
rect 8668 3596 8720 3602
rect 8668 3538 8720 3544
rect 8864 3466 8892 5102
rect 9048 4729 9076 5102
rect 9034 4720 9090 4729
rect 9034 4655 9090 4664
rect 8852 3460 8904 3466
rect 8852 3402 8904 3408
rect 8944 3392 8996 3398
rect 8944 3334 8996 3340
rect 9312 3392 9364 3398
rect 9312 3334 9364 3340
rect 8956 3126 8984 3334
rect 8944 3120 8996 3126
rect 8944 3062 8996 3068
rect 9036 3052 9088 3058
rect 9036 2994 9088 3000
rect 6092 2440 6144 2446
rect 6092 2382 6144 2388
rect 6276 2440 6328 2446
rect 6276 2382 6328 2388
rect 7840 2440 7892 2446
rect 7840 2382 7892 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 4068 2372 4120 2378
rect 4068 2314 4120 2320
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 3737 2204 4045 2213
rect 3737 2202 3743 2204
rect 3799 2202 3823 2204
rect 3879 2202 3903 2204
rect 3959 2202 3983 2204
rect 4039 2202 4045 2204
rect 3799 2150 3801 2202
rect 3981 2150 3983 2202
rect 3737 2148 3743 2150
rect 3799 2148 3823 2150
rect 3879 2148 3903 2150
rect 3959 2148 3983 2150
rect 4039 2148 4045 2150
rect 3737 2139 4045 2148
rect 4080 1170 4108 2314
rect 6460 2304 6512 2310
rect 6460 2246 6512 2252
rect 7104 2304 7156 2310
rect 7104 2246 7156 2252
rect 3896 1142 4108 1170
rect 3896 800 3924 1142
rect 6472 800 6500 2246
rect 7116 800 7144 2246
rect 7992 2204 8300 2213
rect 7992 2202 7998 2204
rect 8054 2202 8078 2204
rect 8134 2202 8158 2204
rect 8214 2202 8238 2204
rect 8294 2202 8300 2204
rect 8054 2150 8056 2202
rect 8236 2150 8238 2202
rect 7992 2148 7998 2150
rect 8054 2148 8078 2150
rect 8134 2148 8158 2150
rect 8214 2148 8238 2150
rect 8294 2148 8300 2150
rect 7992 2139 8300 2148
rect 8404 800 8432 2314
rect 9048 800 9076 2994
rect 9324 2446 9352 3334
rect 9416 2854 9444 8434
rect 10060 8430 10088 8910
rect 10244 8566 10272 8910
rect 10232 8560 10284 8566
rect 10232 8502 10284 8508
rect 10244 8430 10272 8502
rect 10048 8424 10100 8430
rect 10048 8366 10100 8372
rect 10232 8424 10284 8430
rect 10232 8366 10284 8372
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9508 6905 9536 8230
rect 10324 7744 10376 7750
rect 10324 7686 10376 7692
rect 10336 7546 10364 7686
rect 10324 7540 10376 7546
rect 10324 7482 10376 7488
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9494 6896 9550 6905
rect 9494 6831 9550 6840
rect 9600 6798 9628 7414
rect 9772 7404 9824 7410
rect 9772 7346 9824 7352
rect 9588 6792 9640 6798
rect 9588 6734 9640 6740
rect 9784 6662 9812 7346
rect 9954 6896 10010 6905
rect 9954 6831 10010 6840
rect 9968 6798 9996 6831
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 9588 6656 9640 6662
rect 9588 6598 9640 6604
rect 9772 6656 9824 6662
rect 9772 6598 9824 6604
rect 9496 5772 9548 5778
rect 9496 5714 9548 5720
rect 9508 4758 9536 5714
rect 9600 5234 9628 6598
rect 9784 6186 9812 6598
rect 9772 6180 9824 6186
rect 9772 6122 9824 6128
rect 9588 5228 9640 5234
rect 9588 5170 9640 5176
rect 9772 5160 9824 5166
rect 9772 5102 9824 5108
rect 10140 5160 10192 5166
rect 10140 5102 10192 5108
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 9496 4752 9548 4758
rect 9496 4694 9548 4700
rect 9692 4486 9720 5034
rect 9784 4690 9812 5102
rect 9772 4684 9824 4690
rect 9772 4626 9824 4632
rect 9864 4684 9916 4690
rect 9864 4626 9916 4632
rect 9680 4480 9732 4486
rect 9680 4422 9732 4428
rect 9784 4146 9812 4626
rect 9876 4282 9904 4626
rect 10152 4622 10180 5102
rect 10244 4690 10272 5102
rect 10336 4706 10364 7482
rect 10428 5370 10456 9318
rect 10520 8838 10548 13382
rect 10600 13320 10652 13326
rect 10600 13262 10652 13268
rect 10692 13320 10744 13326
rect 10692 13262 10744 13268
rect 10612 12442 10640 13262
rect 10600 12436 10652 12442
rect 10600 12378 10652 12384
rect 10704 12306 10732 13262
rect 10876 12844 10928 12850
rect 10876 12786 10928 12792
rect 10692 12300 10744 12306
rect 10692 12242 10744 12248
rect 10782 10840 10838 10849
rect 10782 10775 10784 10784
rect 10836 10775 10838 10784
rect 10784 10746 10836 10752
rect 10888 10062 10916 12786
rect 10980 10742 11008 13926
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11164 11642 11192 13806
rect 11348 13394 11376 14418
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11244 12844 11296 12850
rect 11244 12786 11296 12792
rect 11256 12238 11284 12786
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11072 11614 11192 11642
rect 10968 10736 11020 10742
rect 10968 10678 11020 10684
rect 10876 10056 10928 10062
rect 10876 9998 10928 10004
rect 10690 9616 10746 9625
rect 10690 9551 10746 9560
rect 10784 9580 10836 9586
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10612 7206 10640 8026
rect 10600 7200 10652 7206
rect 10600 7142 10652 7148
rect 10612 7002 10640 7142
rect 10600 6996 10652 7002
rect 10600 6938 10652 6944
rect 10508 6928 10560 6934
rect 10508 6870 10560 6876
rect 10520 6798 10548 6870
rect 10508 6792 10560 6798
rect 10508 6734 10560 6740
rect 10416 5364 10468 5370
rect 10416 5306 10468 5312
rect 10416 5160 10468 5166
rect 10416 5102 10468 5108
rect 10428 4826 10456 5102
rect 10416 4820 10468 4826
rect 10416 4762 10468 4768
rect 10336 4690 10456 4706
rect 10232 4684 10284 4690
rect 10336 4684 10468 4690
rect 10336 4678 10416 4684
rect 10232 4626 10284 4632
rect 10416 4626 10468 4632
rect 10140 4616 10192 4622
rect 10140 4558 10192 4564
rect 9864 4276 9916 4282
rect 9864 4218 9916 4224
rect 9772 4140 9824 4146
rect 9772 4082 9824 4088
rect 9956 4140 10008 4146
rect 9956 4082 10008 4088
rect 9680 4072 9732 4078
rect 9680 4014 9732 4020
rect 9692 3194 9720 4014
rect 9968 3194 9996 4082
rect 10152 4078 10180 4558
rect 10416 4480 10468 4486
rect 10416 4422 10468 4428
rect 10140 4072 10192 4078
rect 10140 4014 10192 4020
rect 10140 3936 10192 3942
rect 10140 3878 10192 3884
rect 10152 3602 10180 3878
rect 10428 3602 10456 4422
rect 10704 3942 10732 9551
rect 10784 9522 10836 9528
rect 10796 9178 10824 9522
rect 11072 9382 11100 11614
rect 11152 11552 11204 11558
rect 11152 11494 11204 11500
rect 11164 10674 11192 11494
rect 11256 10996 11284 12174
rect 11348 11150 11376 13330
rect 11440 12458 11468 16918
rect 11587 16892 11895 16901
rect 11587 16890 11593 16892
rect 11649 16890 11673 16892
rect 11729 16890 11753 16892
rect 11809 16890 11833 16892
rect 11889 16890 11895 16892
rect 11649 16838 11651 16890
rect 11831 16838 11833 16890
rect 11587 16836 11593 16838
rect 11649 16836 11673 16838
rect 11729 16836 11753 16838
rect 11809 16836 11833 16838
rect 11889 16836 11895 16838
rect 11587 16827 11895 16836
rect 11992 16658 12020 18362
rect 12636 18086 12664 18702
rect 12900 18624 12952 18630
rect 12900 18566 12952 18572
rect 12624 18080 12676 18086
rect 12624 18022 12676 18028
rect 12440 17808 12492 17814
rect 12440 17750 12492 17756
rect 12452 17678 12480 17750
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12247 17436 12555 17445
rect 12247 17434 12253 17436
rect 12309 17434 12333 17436
rect 12389 17434 12413 17436
rect 12469 17434 12493 17436
rect 12549 17434 12555 17436
rect 12309 17382 12311 17434
rect 12491 17382 12493 17434
rect 12247 17380 12253 17382
rect 12309 17380 12333 17382
rect 12389 17380 12413 17382
rect 12469 17380 12493 17382
rect 12549 17380 12555 17382
rect 12247 17371 12555 17380
rect 12636 17354 12664 18022
rect 12912 17678 12940 18566
rect 13096 18426 13124 18702
rect 13636 18624 13688 18630
rect 13636 18566 13688 18572
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13648 18358 13676 18566
rect 13636 18352 13688 18358
rect 13636 18294 13688 18300
rect 13832 17882 13860 18702
rect 14096 18692 14148 18698
rect 14096 18634 14148 18640
rect 13820 17876 13872 17882
rect 13820 17818 13872 17824
rect 13176 17740 13228 17746
rect 13176 17682 13228 17688
rect 12900 17672 12952 17678
rect 12900 17614 12952 17620
rect 12636 17326 12848 17354
rect 11980 16652 12032 16658
rect 11980 16594 12032 16600
rect 12532 16652 12584 16658
rect 12584 16612 12756 16640
rect 12532 16594 12584 16600
rect 11612 16584 11664 16590
rect 11612 16526 11664 16532
rect 11520 16516 11572 16522
rect 11520 16458 11572 16464
rect 11532 16250 11560 16458
rect 11624 16250 11652 16526
rect 11520 16244 11572 16250
rect 11520 16186 11572 16192
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11888 16108 11940 16114
rect 11992 16096 12020 16594
rect 12072 16584 12124 16590
rect 12072 16526 12124 16532
rect 12084 16454 12112 16526
rect 12072 16448 12124 16454
rect 12072 16390 12124 16396
rect 12084 16114 12112 16390
rect 12247 16348 12555 16357
rect 12247 16346 12253 16348
rect 12309 16346 12333 16348
rect 12389 16346 12413 16348
rect 12469 16346 12493 16348
rect 12549 16346 12555 16348
rect 12309 16294 12311 16346
rect 12491 16294 12493 16346
rect 12247 16292 12253 16294
rect 12309 16292 12333 16294
rect 12389 16292 12413 16294
rect 12469 16292 12493 16294
rect 12549 16292 12555 16294
rect 12247 16283 12555 16292
rect 11940 16068 12020 16096
rect 12072 16108 12124 16114
rect 11888 16050 11940 16056
rect 12072 16050 12124 16056
rect 12728 15994 12756 16612
rect 12820 16590 12848 17326
rect 13188 17134 13216 17682
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 12900 16652 12952 16658
rect 12900 16594 12952 16600
rect 13084 16652 13136 16658
rect 13084 16594 13136 16600
rect 12808 16584 12860 16590
rect 12808 16526 12860 16532
rect 12820 16114 12848 16526
rect 12912 16114 12940 16594
rect 12808 16108 12860 16114
rect 12808 16050 12860 16056
rect 12900 16108 12952 16114
rect 12900 16050 12952 16056
rect 12532 15972 12584 15978
rect 12728 15966 12848 15994
rect 12532 15914 12584 15920
rect 11587 15804 11895 15813
rect 11587 15802 11593 15804
rect 11649 15802 11673 15804
rect 11729 15802 11753 15804
rect 11809 15802 11833 15804
rect 11889 15802 11895 15804
rect 11649 15750 11651 15802
rect 11831 15750 11833 15802
rect 11587 15748 11593 15750
rect 11649 15748 11673 15750
rect 11729 15748 11753 15750
rect 11809 15748 11833 15750
rect 11889 15748 11895 15750
rect 11587 15739 11895 15748
rect 12544 15570 12572 15914
rect 12532 15564 12584 15570
rect 12532 15506 12584 15512
rect 12716 15496 12768 15502
rect 12716 15438 12768 15444
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12247 15260 12555 15269
rect 12247 15258 12253 15260
rect 12309 15258 12333 15260
rect 12389 15258 12413 15260
rect 12469 15258 12493 15260
rect 12549 15258 12555 15260
rect 12309 15206 12311 15258
rect 12491 15206 12493 15258
rect 12247 15204 12253 15206
rect 12309 15204 12333 15206
rect 12389 15204 12413 15206
rect 12469 15204 12493 15206
rect 12549 15204 12555 15206
rect 12247 15195 12555 15204
rect 12164 14816 12216 14822
rect 12164 14758 12216 14764
rect 11587 14716 11895 14725
rect 11587 14714 11593 14716
rect 11649 14714 11673 14716
rect 11729 14714 11753 14716
rect 11809 14714 11833 14716
rect 11889 14714 11895 14716
rect 11649 14662 11651 14714
rect 11831 14662 11833 14714
rect 11587 14660 11593 14662
rect 11649 14660 11673 14662
rect 11729 14660 11753 14662
rect 11809 14660 11833 14662
rect 11889 14660 11895 14662
rect 11587 14651 11895 14660
rect 12072 14272 12124 14278
rect 12072 14214 12124 14220
rect 12084 14006 12112 14214
rect 12176 14006 12204 14758
rect 12247 14172 12555 14181
rect 12247 14170 12253 14172
rect 12309 14170 12333 14172
rect 12389 14170 12413 14172
rect 12469 14170 12493 14172
rect 12549 14170 12555 14172
rect 12309 14118 12311 14170
rect 12491 14118 12493 14170
rect 12247 14116 12253 14118
rect 12309 14116 12333 14118
rect 12389 14116 12413 14118
rect 12469 14116 12493 14118
rect 12549 14116 12555 14118
rect 12247 14107 12555 14116
rect 12636 14074 12664 15302
rect 12728 15065 12756 15438
rect 12820 15434 12848 15966
rect 13096 15502 13124 16594
rect 13084 15496 13136 15502
rect 13084 15438 13136 15444
rect 12808 15428 12860 15434
rect 12808 15370 12860 15376
rect 12714 15056 12770 15065
rect 12714 14991 12770 15000
rect 12728 14958 12756 14991
rect 12716 14952 12768 14958
rect 12716 14894 12768 14900
rect 12624 14068 12676 14074
rect 12624 14010 12676 14016
rect 12072 14000 12124 14006
rect 12072 13942 12124 13948
rect 12164 14000 12216 14006
rect 12164 13942 12216 13948
rect 11587 13628 11895 13637
rect 11587 13626 11593 13628
rect 11649 13626 11673 13628
rect 11729 13626 11753 13628
rect 11809 13626 11833 13628
rect 11889 13626 11895 13628
rect 11649 13574 11651 13626
rect 11831 13574 11833 13626
rect 11587 13572 11593 13574
rect 11649 13572 11673 13574
rect 11729 13572 11753 13574
rect 11809 13572 11833 13574
rect 11889 13572 11895 13574
rect 11587 13563 11895 13572
rect 12084 12986 12112 13942
rect 12624 13932 12676 13938
rect 12624 13874 12676 13880
rect 12440 13728 12492 13734
rect 12440 13670 12492 13676
rect 12452 13326 12480 13670
rect 12440 13320 12492 13326
rect 12440 13262 12492 13268
rect 12247 13084 12555 13093
rect 12247 13082 12253 13084
rect 12309 13082 12333 13084
rect 12389 13082 12413 13084
rect 12469 13082 12493 13084
rect 12549 13082 12555 13084
rect 12309 13030 12311 13082
rect 12491 13030 12493 13082
rect 12247 13028 12253 13030
rect 12309 13028 12333 13030
rect 12389 13028 12413 13030
rect 12469 13028 12493 13030
rect 12549 13028 12555 13030
rect 12247 13019 12555 13028
rect 12636 12986 12664 13874
rect 12992 13388 13044 13394
rect 12992 13330 13044 13336
rect 12808 13184 12860 13190
rect 12808 13126 12860 13132
rect 12072 12980 12124 12986
rect 12072 12922 12124 12928
rect 12624 12980 12676 12986
rect 12624 12922 12676 12928
rect 12820 12918 12848 13126
rect 12808 12912 12860 12918
rect 12808 12854 12860 12860
rect 12440 12844 12492 12850
rect 12440 12786 12492 12792
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12072 12776 12124 12782
rect 12124 12736 12204 12764
rect 12072 12718 12124 12724
rect 11587 12540 11895 12549
rect 11587 12538 11593 12540
rect 11649 12538 11673 12540
rect 11729 12538 11753 12540
rect 11809 12538 11833 12540
rect 11889 12538 11895 12540
rect 11649 12486 11651 12538
rect 11831 12486 11833 12538
rect 11587 12484 11593 12486
rect 11649 12484 11673 12486
rect 11729 12484 11753 12486
rect 11809 12484 11833 12486
rect 11889 12484 11895 12486
rect 11587 12475 11895 12484
rect 11440 12430 11560 12458
rect 11428 11756 11480 11762
rect 11428 11698 11480 11704
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11336 11008 11388 11014
rect 11256 10968 11336 10996
rect 11336 10950 11388 10956
rect 11152 10668 11204 10674
rect 11152 10610 11204 10616
rect 11348 10130 11376 10950
rect 11440 10810 11468 11698
rect 11532 11506 11560 12430
rect 12176 11778 12204 12736
rect 12452 12238 12480 12786
rect 12624 12640 12676 12646
rect 12624 12582 12676 12588
rect 12440 12232 12492 12238
rect 12440 12174 12492 12180
rect 12636 12102 12664 12582
rect 12728 12170 12756 12786
rect 13004 12646 13032 13330
rect 12992 12640 13044 12646
rect 12992 12582 13044 12588
rect 13004 12442 13032 12582
rect 12992 12436 13044 12442
rect 12992 12378 13044 12384
rect 12808 12232 12860 12238
rect 12808 12174 12860 12180
rect 12716 12164 12768 12170
rect 12716 12106 12768 12112
rect 12624 12096 12676 12102
rect 12624 12038 12676 12044
rect 12247 11996 12555 12005
rect 12247 11994 12253 11996
rect 12309 11994 12333 11996
rect 12389 11994 12413 11996
rect 12469 11994 12493 11996
rect 12549 11994 12555 11996
rect 12309 11942 12311 11994
rect 12491 11942 12493 11994
rect 12247 11940 12253 11942
rect 12309 11940 12333 11942
rect 12389 11940 12413 11942
rect 12469 11940 12493 11942
rect 12549 11940 12555 11942
rect 12247 11931 12555 11940
rect 11523 11478 11560 11506
rect 11992 11750 12204 11778
rect 11523 11370 11551 11478
rect 11587 11452 11895 11461
rect 11587 11450 11593 11452
rect 11649 11450 11673 11452
rect 11729 11450 11753 11452
rect 11809 11450 11833 11452
rect 11889 11450 11895 11452
rect 11649 11398 11651 11450
rect 11831 11398 11833 11450
rect 11587 11396 11593 11398
rect 11649 11396 11673 11398
rect 11729 11396 11753 11398
rect 11809 11396 11833 11398
rect 11889 11396 11895 11398
rect 11587 11387 11895 11396
rect 11523 11342 11560 11370
rect 11428 10804 11480 10810
rect 11428 10746 11480 10752
rect 11532 10418 11560 11342
rect 11992 10674 12020 11750
rect 12256 11552 12308 11558
rect 12256 11494 12308 11500
rect 12624 11552 12676 11558
rect 12624 11494 12676 11500
rect 12268 11150 12296 11494
rect 12636 11150 12664 11494
rect 12256 11144 12308 11150
rect 12256 11086 12308 11092
rect 12624 11144 12676 11150
rect 12624 11086 12676 11092
rect 12072 11076 12124 11082
rect 12072 11018 12124 11024
rect 12084 10810 12112 11018
rect 12636 11014 12664 11086
rect 12624 11008 12676 11014
rect 12624 10950 12676 10956
rect 12247 10908 12555 10917
rect 12247 10906 12253 10908
rect 12309 10906 12333 10908
rect 12389 10906 12413 10908
rect 12469 10906 12493 10908
rect 12549 10906 12555 10908
rect 12309 10854 12311 10906
rect 12491 10854 12493 10906
rect 12247 10852 12253 10854
rect 12309 10852 12333 10854
rect 12389 10852 12413 10854
rect 12469 10852 12493 10854
rect 12549 10852 12555 10854
rect 12247 10843 12555 10852
rect 12072 10804 12124 10810
rect 12072 10746 12124 10752
rect 11980 10668 12032 10674
rect 11980 10610 12032 10616
rect 12256 10600 12308 10606
rect 12256 10542 12308 10548
rect 11523 10390 11560 10418
rect 11523 10282 11551 10390
rect 11587 10364 11895 10373
rect 11587 10362 11593 10364
rect 11649 10362 11673 10364
rect 11729 10362 11753 10364
rect 11809 10362 11833 10364
rect 11889 10362 11895 10364
rect 11649 10310 11651 10362
rect 11831 10310 11833 10362
rect 11587 10308 11593 10310
rect 11649 10308 11673 10310
rect 11729 10308 11753 10310
rect 11809 10308 11833 10310
rect 11889 10308 11895 10310
rect 11587 10299 11895 10308
rect 11523 10254 11560 10282
rect 11532 10248 11560 10254
rect 11532 10220 11928 10248
rect 11336 10124 11388 10130
rect 11336 10066 11388 10072
rect 11612 9988 11664 9994
rect 11612 9930 11664 9936
rect 11704 9988 11756 9994
rect 11704 9930 11756 9936
rect 11428 9580 11480 9586
rect 11428 9522 11480 9528
rect 11244 9512 11296 9518
rect 11244 9454 11296 9460
rect 11060 9376 11112 9382
rect 11060 9318 11112 9324
rect 10784 9172 10836 9178
rect 10784 9114 10836 9120
rect 10876 8832 10928 8838
rect 10876 8774 10928 8780
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 10784 8356 10836 8362
rect 10888 8344 10916 8774
rect 11164 8430 11192 8774
rect 11152 8424 11204 8430
rect 11256 8401 11284 9454
rect 11440 9178 11468 9522
rect 11624 9450 11652 9930
rect 11716 9625 11744 9930
rect 11702 9616 11758 9625
rect 11702 9551 11758 9560
rect 11900 9518 11928 10220
rect 12268 9908 12296 10542
rect 12636 10470 12664 10950
rect 12728 10674 12756 12106
rect 12820 11762 12848 12174
rect 12808 11756 12860 11762
rect 12808 11698 12860 11704
rect 12820 11286 12848 11698
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 13096 11354 13124 11562
rect 13084 11348 13136 11354
rect 13084 11290 13136 11296
rect 12808 11280 12860 11286
rect 12808 11222 12860 11228
rect 12716 10668 12768 10674
rect 12716 10610 12768 10616
rect 13084 10668 13136 10674
rect 13084 10610 13136 10616
rect 12624 10464 12676 10470
rect 12624 10406 12676 10412
rect 12624 10260 12676 10266
rect 12624 10202 12676 10208
rect 12176 9880 12296 9908
rect 11980 9580 12032 9586
rect 11980 9522 12032 9528
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11612 9444 11664 9450
rect 11612 9386 11664 9392
rect 11587 9276 11895 9285
rect 11587 9274 11593 9276
rect 11649 9274 11673 9276
rect 11729 9274 11753 9276
rect 11809 9274 11833 9276
rect 11889 9274 11895 9276
rect 11649 9222 11651 9274
rect 11831 9222 11833 9274
rect 11587 9220 11593 9222
rect 11649 9220 11673 9222
rect 11729 9220 11753 9222
rect 11809 9220 11833 9222
rect 11889 9220 11895 9222
rect 11587 9211 11895 9220
rect 11428 9172 11480 9178
rect 11428 9114 11480 9120
rect 11888 8832 11940 8838
rect 11888 8774 11940 8780
rect 11900 8514 11928 8774
rect 11992 8634 12020 9522
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 8906 12112 9318
rect 12072 8900 12124 8906
rect 12072 8842 12124 8848
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 11900 8486 12020 8514
rect 11152 8366 11204 8372
rect 11242 8392 11298 8401
rect 10836 8316 10916 8344
rect 11242 8327 11298 8336
rect 10784 8298 10836 8304
rect 10784 6724 10836 6730
rect 10784 6666 10836 6672
rect 10796 6458 10824 6666
rect 10784 6452 10836 6458
rect 10784 6394 10836 6400
rect 10692 3936 10744 3942
rect 10692 3878 10744 3884
rect 10600 3664 10652 3670
rect 10600 3606 10652 3612
rect 10140 3596 10192 3602
rect 10140 3538 10192 3544
rect 10416 3596 10468 3602
rect 10416 3538 10468 3544
rect 9680 3188 9732 3194
rect 9680 3130 9732 3136
rect 9956 3188 10008 3194
rect 9956 3130 10008 3136
rect 10152 2961 10180 3538
rect 10138 2952 10194 2961
rect 10138 2887 10194 2896
rect 9404 2848 9456 2854
rect 9404 2790 9456 2796
rect 10428 2650 10456 3538
rect 10612 3058 10640 3606
rect 10600 3052 10652 3058
rect 10600 2994 10652 3000
rect 10416 2644 10468 2650
rect 10416 2586 10468 2592
rect 10888 2514 10916 8316
rect 11060 7744 11112 7750
rect 11060 7686 11112 7692
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 10980 5710 11008 6598
rect 11072 6390 11100 7686
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 11164 6322 11192 7142
rect 11152 6316 11204 6322
rect 11152 6258 11204 6264
rect 11256 5794 11284 8327
rect 11587 8188 11895 8197
rect 11587 8186 11593 8188
rect 11649 8186 11673 8188
rect 11729 8186 11753 8188
rect 11809 8186 11833 8188
rect 11889 8186 11895 8188
rect 11649 8134 11651 8186
rect 11831 8134 11833 8186
rect 11587 8132 11593 8134
rect 11649 8132 11673 8134
rect 11729 8132 11753 8134
rect 11809 8132 11833 8134
rect 11889 8132 11895 8134
rect 11587 8123 11895 8132
rect 11992 8072 12020 8486
rect 12176 8430 12204 9880
rect 12247 9820 12555 9829
rect 12247 9818 12253 9820
rect 12309 9818 12333 9820
rect 12389 9818 12413 9820
rect 12469 9818 12493 9820
rect 12549 9818 12555 9820
rect 12309 9766 12311 9818
rect 12491 9766 12493 9818
rect 12247 9764 12253 9766
rect 12309 9764 12333 9766
rect 12389 9764 12413 9766
rect 12469 9764 12493 9766
rect 12549 9764 12555 9766
rect 12247 9755 12555 9764
rect 12636 9178 12664 10202
rect 12624 9172 12676 9178
rect 12624 9114 12676 9120
rect 12624 8900 12676 8906
rect 12624 8842 12676 8848
rect 12247 8732 12555 8741
rect 12247 8730 12253 8732
rect 12309 8730 12333 8732
rect 12389 8730 12413 8732
rect 12469 8730 12493 8732
rect 12549 8730 12555 8732
rect 12309 8678 12311 8730
rect 12491 8678 12493 8730
rect 12247 8676 12253 8678
rect 12309 8676 12333 8678
rect 12389 8676 12413 8678
rect 12469 8676 12493 8678
rect 12549 8676 12555 8678
rect 12247 8667 12555 8676
rect 12164 8424 12216 8430
rect 12164 8366 12216 8372
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 11900 8044 12020 8072
rect 11900 7290 11928 8044
rect 12084 7478 12112 8230
rect 12532 7880 12584 7886
rect 12530 7848 12532 7857
rect 12584 7848 12586 7857
rect 12530 7783 12586 7792
rect 12247 7644 12555 7653
rect 12247 7642 12253 7644
rect 12309 7642 12333 7644
rect 12389 7642 12413 7644
rect 12469 7642 12493 7644
rect 12549 7642 12555 7644
rect 12309 7590 12311 7642
rect 12491 7590 12493 7642
rect 12247 7588 12253 7590
rect 12309 7588 12333 7590
rect 12389 7588 12413 7590
rect 12469 7588 12493 7590
rect 12549 7588 12555 7590
rect 12247 7579 12555 7588
rect 12072 7472 12124 7478
rect 11978 7440 12034 7449
rect 12072 7414 12124 7420
rect 11978 7375 11980 7384
rect 12032 7375 12034 7384
rect 12164 7404 12216 7410
rect 11980 7346 12032 7352
rect 12164 7346 12216 7352
rect 12348 7404 12400 7410
rect 12348 7346 12400 7352
rect 12532 7404 12584 7410
rect 12532 7346 12584 7352
rect 11900 7262 12112 7290
rect 12176 7274 12204 7346
rect 11587 7100 11895 7109
rect 11587 7098 11593 7100
rect 11649 7098 11673 7100
rect 11729 7098 11753 7100
rect 11809 7098 11833 7100
rect 11889 7098 11895 7100
rect 11649 7046 11651 7098
rect 11831 7046 11833 7098
rect 11587 7044 11593 7046
rect 11649 7044 11673 7046
rect 11729 7044 11753 7046
rect 11809 7044 11833 7046
rect 11889 7044 11895 7046
rect 11587 7035 11895 7044
rect 11888 6792 11940 6798
rect 11886 6760 11888 6769
rect 11940 6760 11942 6769
rect 11886 6695 11942 6704
rect 11900 6361 11928 6695
rect 11886 6352 11942 6361
rect 11886 6287 11942 6296
rect 11336 6248 11388 6254
rect 11336 6190 11388 6196
rect 11348 5914 11376 6190
rect 11428 6112 11480 6118
rect 11428 6054 11480 6060
rect 11336 5908 11388 5914
rect 11336 5850 11388 5856
rect 11060 5772 11112 5778
rect 11060 5714 11112 5720
rect 11152 5772 11204 5778
rect 11256 5766 11376 5794
rect 11152 5714 11204 5720
rect 10968 5704 11020 5710
rect 10968 5646 11020 5652
rect 11072 5370 11100 5714
rect 10968 5364 11020 5370
rect 10968 5306 11020 5312
rect 11060 5364 11112 5370
rect 11060 5306 11112 5312
rect 10980 4146 11008 5306
rect 11164 4826 11192 5714
rect 11244 5704 11296 5710
rect 11242 5672 11244 5681
rect 11296 5672 11298 5681
rect 11242 5607 11298 5616
rect 11348 5114 11376 5766
rect 11440 5710 11468 6054
rect 11587 6012 11895 6021
rect 11587 6010 11593 6012
rect 11649 6010 11673 6012
rect 11729 6010 11753 6012
rect 11809 6010 11833 6012
rect 11889 6010 11895 6012
rect 11649 5958 11651 6010
rect 11831 5958 11833 6010
rect 11587 5956 11593 5958
rect 11649 5956 11673 5958
rect 11729 5956 11753 5958
rect 11809 5956 11833 5958
rect 11889 5956 11895 5958
rect 11587 5947 11895 5956
rect 11428 5704 11480 5710
rect 11428 5646 11480 5652
rect 11428 5228 11480 5234
rect 11428 5170 11480 5176
rect 11256 5086 11376 5114
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 10968 4140 11020 4146
rect 10968 4082 11020 4088
rect 11256 4010 11284 5086
rect 11336 5024 11388 5030
rect 11336 4966 11388 4972
rect 11348 4554 11376 4966
rect 11336 4548 11388 4554
rect 11336 4490 11388 4496
rect 11440 4282 11468 5170
rect 11587 4924 11895 4933
rect 11587 4922 11593 4924
rect 11649 4922 11673 4924
rect 11729 4922 11753 4924
rect 11809 4922 11833 4924
rect 11889 4922 11895 4924
rect 11649 4870 11651 4922
rect 11831 4870 11833 4922
rect 11587 4868 11593 4870
rect 11649 4868 11673 4870
rect 11729 4868 11753 4870
rect 11809 4868 11833 4870
rect 11889 4868 11895 4870
rect 11587 4859 11895 4868
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11244 4004 11296 4010
rect 11244 3946 11296 3952
rect 10968 3936 11020 3942
rect 10968 3878 11020 3884
rect 10980 3534 11008 3878
rect 11256 3602 11284 3946
rect 11980 3936 12032 3942
rect 11980 3878 12032 3884
rect 11587 3836 11895 3845
rect 11587 3834 11593 3836
rect 11649 3834 11673 3836
rect 11729 3834 11753 3836
rect 11809 3834 11833 3836
rect 11889 3834 11895 3836
rect 11649 3782 11651 3834
rect 11831 3782 11833 3834
rect 11587 3780 11593 3782
rect 11649 3780 11673 3782
rect 11729 3780 11753 3782
rect 11809 3780 11833 3782
rect 11889 3780 11895 3782
rect 11587 3771 11895 3780
rect 11244 3596 11296 3602
rect 11244 3538 11296 3544
rect 10968 3528 11020 3534
rect 10968 3470 11020 3476
rect 11992 3058 12020 3878
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 11587 2748 11895 2757
rect 11587 2746 11593 2748
rect 11649 2746 11673 2748
rect 11729 2746 11753 2748
rect 11809 2746 11833 2748
rect 11889 2746 11895 2748
rect 11649 2694 11651 2746
rect 11831 2694 11833 2746
rect 11587 2692 11593 2694
rect 11649 2692 11673 2694
rect 11729 2692 11753 2694
rect 11809 2692 11833 2694
rect 11889 2692 11895 2694
rect 11587 2683 11895 2692
rect 11612 2576 11664 2582
rect 11612 2518 11664 2524
rect 10876 2508 10928 2514
rect 10876 2450 10928 2456
rect 9312 2440 9364 2446
rect 9312 2382 9364 2388
rect 10324 2440 10376 2446
rect 10324 2382 10376 2388
rect 9680 2372 9732 2378
rect 9680 2314 9732 2320
rect 9692 800 9720 2314
rect 10336 800 10364 2382
rect 10968 2304 11020 2310
rect 10968 2246 11020 2252
rect 10980 800 11008 2246
rect 11624 800 11652 2518
rect 12084 2514 12112 7262
rect 12164 7268 12216 7274
rect 12164 7210 12216 7216
rect 12176 6866 12204 7210
rect 12360 7002 12388 7346
rect 12544 7206 12572 7346
rect 12532 7200 12584 7206
rect 12532 7142 12584 7148
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12164 6860 12216 6866
rect 12164 6802 12216 6808
rect 12636 6662 12664 8842
rect 12728 8090 12756 10610
rect 12806 10296 12862 10305
rect 12806 10231 12808 10240
rect 12860 10231 12862 10240
rect 12808 10202 12860 10208
rect 12820 9654 12848 10202
rect 12808 9648 12860 9654
rect 12808 9590 12860 9596
rect 12716 8084 12768 8090
rect 12716 8026 12768 8032
rect 12820 7970 12848 9590
rect 12992 9036 13044 9042
rect 12992 8978 13044 8984
rect 12900 8560 12952 8566
rect 12900 8502 12952 8508
rect 12728 7942 12848 7970
rect 12728 7750 12756 7942
rect 12808 7812 12860 7818
rect 12808 7754 12860 7760
rect 12716 7744 12768 7750
rect 12716 7686 12768 7692
rect 12716 7540 12768 7546
rect 12716 7482 12768 7488
rect 12728 7410 12756 7482
rect 12820 7410 12848 7754
rect 12716 7404 12768 7410
rect 12716 7346 12768 7352
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12912 7206 12940 8502
rect 13004 8090 13032 8978
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 13004 7478 13032 7686
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 13096 7410 13124 10610
rect 13188 10062 13216 17070
rect 13268 15904 13320 15910
rect 13268 15846 13320 15852
rect 13280 13938 13308 15846
rect 13912 15496 13964 15502
rect 13912 15438 13964 15444
rect 13728 15428 13780 15434
rect 13728 15370 13780 15376
rect 13740 15178 13768 15370
rect 13740 15150 13860 15178
rect 13924 15162 13952 15438
rect 13832 14793 13860 15150
rect 13912 15156 13964 15162
rect 13912 15098 13964 15104
rect 13924 15026 13952 15098
rect 13912 15020 13964 15026
rect 13912 14962 13964 14968
rect 13818 14784 13874 14793
rect 13818 14719 13874 14728
rect 14108 14618 14136 18634
rect 16502 18524 16810 18533
rect 16502 18522 16508 18524
rect 16564 18522 16588 18524
rect 16644 18522 16668 18524
rect 16724 18522 16748 18524
rect 16804 18522 16810 18524
rect 16564 18470 16566 18522
rect 16746 18470 16748 18522
rect 16502 18468 16508 18470
rect 16564 18468 16588 18470
rect 16644 18468 16668 18470
rect 16724 18468 16748 18470
rect 16804 18468 16810 18470
rect 16502 18459 16810 18468
rect 15660 18284 15712 18290
rect 15660 18226 15712 18232
rect 15016 18148 15068 18154
rect 15016 18090 15068 18096
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14752 17610 14780 18022
rect 14924 17672 14976 17678
rect 14924 17614 14976 17620
rect 14740 17604 14792 17610
rect 14740 17546 14792 17552
rect 14464 17536 14516 17542
rect 14464 17478 14516 17484
rect 14556 17536 14608 17542
rect 14556 17478 14608 17484
rect 14476 17338 14504 17478
rect 14568 17338 14596 17478
rect 14464 17332 14516 17338
rect 14464 17274 14516 17280
rect 14556 17332 14608 17338
rect 14556 17274 14608 17280
rect 14464 16652 14516 16658
rect 14464 16594 14516 16600
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 13452 14408 13504 14414
rect 13452 14350 13504 14356
rect 13268 13932 13320 13938
rect 13268 13874 13320 13880
rect 13268 13252 13320 13258
rect 13268 13194 13320 13200
rect 13360 13252 13412 13258
rect 13360 13194 13412 13200
rect 13280 12850 13308 13194
rect 13372 12850 13400 13194
rect 13268 12844 13320 12850
rect 13268 12786 13320 12792
rect 13360 12844 13412 12850
rect 13360 12786 13412 12792
rect 13280 10810 13308 12786
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13372 10690 13400 12786
rect 13464 10810 13492 14350
rect 13728 14340 13780 14346
rect 13728 14282 13780 14288
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13556 12918 13584 14010
rect 13740 13841 13768 14282
rect 14292 13938 14320 15302
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14384 14793 14412 14826
rect 14370 14784 14426 14793
rect 14370 14719 14426 14728
rect 14476 14618 14504 16594
rect 14936 16182 14964 17614
rect 14924 16176 14976 16182
rect 14924 16118 14976 16124
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14752 15502 14780 15846
rect 15028 15502 15056 18090
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15396 17678 15424 18022
rect 15384 17672 15436 17678
rect 15384 17614 15436 17620
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15108 17264 15160 17270
rect 15108 17206 15160 17212
rect 14740 15496 14792 15502
rect 14740 15438 14792 15444
rect 14832 15496 14884 15502
rect 14832 15438 14884 15444
rect 15016 15496 15068 15502
rect 15016 15438 15068 15444
rect 14844 15162 14872 15438
rect 14832 15156 14884 15162
rect 14832 15098 14884 15104
rect 15028 15026 15056 15438
rect 15016 15020 15068 15026
rect 15016 14962 15068 14968
rect 15120 14822 15148 17206
rect 15580 16658 15608 17614
rect 15672 17338 15700 18226
rect 15842 17980 16150 17989
rect 15842 17978 15848 17980
rect 15904 17978 15928 17980
rect 15984 17978 16008 17980
rect 16064 17978 16088 17980
rect 16144 17978 16150 17980
rect 15904 17926 15906 17978
rect 16086 17926 16088 17978
rect 15842 17924 15848 17926
rect 15904 17924 15928 17926
rect 15984 17924 16008 17926
rect 16064 17924 16088 17926
rect 16144 17924 16150 17926
rect 15842 17915 16150 17924
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 15660 17332 15712 17338
rect 15660 17274 15712 17280
rect 15842 16892 16150 16901
rect 15842 16890 15848 16892
rect 15904 16890 15928 16892
rect 15984 16890 16008 16892
rect 16064 16890 16088 16892
rect 16144 16890 16150 16892
rect 15904 16838 15906 16890
rect 16086 16838 16088 16890
rect 15842 16836 15848 16838
rect 15904 16836 15928 16838
rect 15984 16836 16008 16838
rect 16064 16836 16088 16838
rect 16144 16836 16150 16838
rect 15842 16827 16150 16836
rect 15568 16652 15620 16658
rect 15568 16594 15620 16600
rect 15292 16584 15344 16590
rect 15292 16526 15344 16532
rect 15304 16250 15332 16526
rect 15292 16244 15344 16250
rect 15292 16186 15344 16192
rect 15200 16108 15252 16114
rect 15200 16050 15252 16056
rect 14740 14816 14792 14822
rect 14740 14758 14792 14764
rect 15108 14816 15160 14822
rect 15108 14758 15160 14764
rect 14752 14618 14780 14758
rect 15212 14618 15240 16050
rect 15580 15570 15608 16594
rect 15660 15972 15712 15978
rect 15660 15914 15712 15920
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 14464 14612 14516 14618
rect 14464 14554 14516 14560
rect 14740 14612 14792 14618
rect 14740 14554 14792 14560
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 14372 14408 14424 14414
rect 14372 14350 14424 14356
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 13726 13832 13782 13841
rect 13782 13790 13860 13818
rect 13726 13767 13782 13776
rect 13832 13326 13860 13790
rect 13820 13320 13872 13326
rect 13820 13262 13872 13268
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13728 12844 13780 12850
rect 13728 12786 13780 12792
rect 13740 12442 13768 12786
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13832 11778 13860 12174
rect 13740 11762 13860 11778
rect 13728 11756 13860 11762
rect 13780 11750 13860 11756
rect 13728 11698 13780 11704
rect 13728 11620 13780 11626
rect 13728 11562 13780 11568
rect 13544 11552 13596 11558
rect 13544 11494 13596 11500
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13280 10674 13400 10690
rect 13556 10674 13584 11494
rect 13268 10668 13400 10674
rect 13320 10662 13400 10668
rect 13544 10668 13596 10674
rect 13268 10610 13320 10616
rect 13544 10610 13596 10616
rect 13176 10056 13228 10062
rect 13176 9998 13228 10004
rect 13280 9722 13308 10610
rect 13740 10062 13768 11562
rect 13360 10056 13412 10062
rect 13358 10024 13360 10033
rect 13452 10056 13504 10062
rect 13412 10024 13414 10033
rect 13452 9998 13504 10004
rect 13728 10056 13780 10062
rect 13728 9998 13780 10004
rect 13358 9959 13414 9968
rect 13464 9722 13492 9998
rect 13268 9716 13320 9722
rect 13268 9658 13320 9664
rect 13452 9716 13504 9722
rect 13452 9658 13504 9664
rect 13176 8832 13228 8838
rect 13176 8774 13228 8780
rect 13188 8634 13216 8774
rect 13176 8628 13228 8634
rect 13176 8570 13228 8576
rect 13176 8492 13228 8498
rect 13176 8434 13228 8440
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 12992 7336 13044 7342
rect 12992 7278 13044 7284
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 13004 7002 13032 7278
rect 12992 6996 13044 7002
rect 12992 6938 13044 6944
rect 12624 6656 12676 6662
rect 12624 6598 12676 6604
rect 12247 6556 12555 6565
rect 12247 6554 12253 6556
rect 12309 6554 12333 6556
rect 12389 6554 12413 6556
rect 12469 6554 12493 6556
rect 12549 6554 12555 6556
rect 12309 6502 12311 6554
rect 12491 6502 12493 6554
rect 12247 6500 12253 6502
rect 12309 6500 12333 6502
rect 12389 6500 12413 6502
rect 12469 6500 12493 6502
rect 12549 6500 12555 6502
rect 12247 6491 12555 6500
rect 12636 6322 12664 6598
rect 12440 6316 12492 6322
rect 12440 6258 12492 6264
rect 12624 6316 12676 6322
rect 12624 6258 12676 6264
rect 12256 6248 12308 6254
rect 12256 6190 12308 6196
rect 12268 5710 12296 6190
rect 12452 5710 12480 6258
rect 12256 5704 12308 5710
rect 12256 5646 12308 5652
rect 12440 5704 12492 5710
rect 12440 5646 12492 5652
rect 12247 5468 12555 5477
rect 12247 5466 12253 5468
rect 12309 5466 12333 5468
rect 12389 5466 12413 5468
rect 12469 5466 12493 5468
rect 12549 5466 12555 5468
rect 12309 5414 12311 5466
rect 12491 5414 12493 5466
rect 12247 5412 12253 5414
rect 12309 5412 12333 5414
rect 12389 5412 12413 5414
rect 12469 5412 12493 5414
rect 12549 5412 12555 5414
rect 12247 5403 12555 5412
rect 12636 4622 12664 6258
rect 13096 6186 13124 7346
rect 13084 6180 13136 6186
rect 13084 6122 13136 6128
rect 12992 5772 13044 5778
rect 12992 5714 13044 5720
rect 12716 5636 12768 5642
rect 12716 5578 12768 5584
rect 12728 5098 12756 5578
rect 12808 5160 12860 5166
rect 12808 5102 12860 5108
rect 12716 5092 12768 5098
rect 12716 5034 12768 5040
rect 12624 4616 12676 4622
rect 12624 4558 12676 4564
rect 12247 4380 12555 4389
rect 12247 4378 12253 4380
rect 12309 4378 12333 4380
rect 12389 4378 12413 4380
rect 12469 4378 12493 4380
rect 12549 4378 12555 4380
rect 12309 4326 12311 4378
rect 12491 4326 12493 4378
rect 12247 4324 12253 4326
rect 12309 4324 12333 4326
rect 12389 4324 12413 4326
rect 12469 4324 12493 4326
rect 12549 4324 12555 4326
rect 12247 4315 12555 4324
rect 12440 4004 12492 4010
rect 12440 3946 12492 3952
rect 12452 3602 12480 3946
rect 12440 3596 12492 3602
rect 12440 3538 12492 3544
rect 12247 3292 12555 3301
rect 12247 3290 12253 3292
rect 12309 3290 12333 3292
rect 12389 3290 12413 3292
rect 12469 3290 12493 3292
rect 12549 3290 12555 3292
rect 12309 3238 12311 3290
rect 12491 3238 12493 3290
rect 12247 3236 12253 3238
rect 12309 3236 12333 3238
rect 12389 3236 12413 3238
rect 12469 3236 12493 3238
rect 12549 3236 12555 3238
rect 12247 3227 12555 3236
rect 12636 3126 12664 4558
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 12728 4282 12756 4422
rect 12716 4276 12768 4282
rect 12716 4218 12768 4224
rect 12820 4146 12848 5102
rect 12716 4140 12768 4146
rect 12716 4082 12768 4088
rect 12808 4140 12860 4146
rect 12808 4082 12860 4088
rect 12728 3670 12756 4082
rect 12716 3664 12768 3670
rect 12716 3606 12768 3612
rect 12820 3194 12848 4082
rect 12808 3188 12860 3194
rect 12808 3130 12860 3136
rect 12624 3120 12676 3126
rect 12624 3062 12676 3068
rect 13004 3040 13032 5714
rect 13188 5234 13216 8434
rect 13280 7410 13308 9658
rect 13360 9172 13412 9178
rect 13360 9114 13412 9120
rect 13372 8498 13400 9114
rect 13636 8900 13688 8906
rect 13636 8842 13688 8848
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13452 8560 13504 8566
rect 13452 8502 13504 8508
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13464 7886 13492 8502
rect 13452 7880 13504 7886
rect 13452 7822 13504 7828
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13464 6730 13492 7822
rect 13556 7546 13584 8774
rect 13648 8362 13676 8842
rect 13740 8566 13768 9998
rect 13832 9926 13860 11750
rect 13924 10810 13952 13874
rect 14384 12986 14412 14350
rect 15476 14272 15528 14278
rect 15476 14214 15528 14220
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 14464 13932 14516 13938
rect 14464 13874 14516 13880
rect 14476 12986 14504 13874
rect 15200 13864 15252 13870
rect 15304 13852 15332 13942
rect 15252 13824 15332 13852
rect 15200 13806 15252 13812
rect 15108 13796 15160 13802
rect 15108 13738 15160 13744
rect 14556 13728 14608 13734
rect 14556 13670 14608 13676
rect 14648 13728 14700 13734
rect 14648 13670 14700 13676
rect 14568 13274 14596 13670
rect 14660 13462 14688 13670
rect 14648 13456 14700 13462
rect 14648 13398 14700 13404
rect 14568 13246 14688 13274
rect 14660 13190 14688 13246
rect 14648 13184 14700 13190
rect 14648 13126 14700 13132
rect 14372 12980 14424 12986
rect 14372 12922 14424 12928
rect 14464 12980 14516 12986
rect 14464 12922 14516 12928
rect 14188 12844 14240 12850
rect 14188 12786 14240 12792
rect 14372 12844 14424 12850
rect 14372 12786 14424 12792
rect 14464 12844 14516 12850
rect 14464 12786 14516 12792
rect 14200 12434 14228 12786
rect 14200 12406 14320 12434
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 14016 11898 14044 12038
rect 14004 11892 14056 11898
rect 14004 11834 14056 11840
rect 14004 11756 14056 11762
rect 14004 11698 14056 11704
rect 13912 10804 13964 10810
rect 13912 10746 13964 10752
rect 13912 10668 13964 10674
rect 13912 10610 13964 10616
rect 13924 10266 13952 10610
rect 13912 10260 13964 10266
rect 13912 10202 13964 10208
rect 14016 10062 14044 11698
rect 14096 11348 14148 11354
rect 14096 11290 14148 11296
rect 14108 10742 14136 11290
rect 14188 11008 14240 11014
rect 14188 10950 14240 10956
rect 14200 10742 14228 10950
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14188 10736 14240 10742
rect 14188 10678 14240 10684
rect 14292 10674 14320 12406
rect 14384 12374 14412 12786
rect 14372 12368 14424 12374
rect 14372 12310 14424 12316
rect 14476 11898 14504 12786
rect 14556 12776 14608 12782
rect 14556 12718 14608 12724
rect 14464 11892 14516 11898
rect 14464 11834 14516 11840
rect 14372 11280 14424 11286
rect 14372 11222 14424 11228
rect 14280 10668 14332 10674
rect 14280 10610 14332 10616
rect 14004 10056 14056 10062
rect 13910 10024 13966 10033
rect 14004 9998 14056 10004
rect 13910 9959 13966 9968
rect 13820 9920 13872 9926
rect 13820 9862 13872 9868
rect 13924 9874 13952 9959
rect 13728 8560 13780 8566
rect 13728 8502 13780 8508
rect 13832 8498 13860 9862
rect 13924 9846 14044 9874
rect 13820 8492 13872 8498
rect 13820 8434 13872 8440
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 13832 8294 13860 8434
rect 13820 8288 13872 8294
rect 13820 8230 13872 8236
rect 13912 8288 13964 8294
rect 13912 8230 13964 8236
rect 13924 7698 13952 8230
rect 14016 7886 14044 9846
rect 14292 8634 14320 10610
rect 14384 8974 14412 11222
rect 14568 10674 14596 12718
rect 14660 11762 14688 13126
rect 14924 12640 14976 12646
rect 14924 12582 14976 12588
rect 14936 12238 14964 12582
rect 15120 12306 15148 13738
rect 15200 13728 15252 13734
rect 15200 13670 15252 13676
rect 15212 12918 15240 13670
rect 15488 13326 15516 14214
rect 15580 13530 15608 15506
rect 15672 14958 15700 15914
rect 15752 15904 15804 15910
rect 15752 15846 15804 15852
rect 15764 15162 15792 15846
rect 15842 15804 16150 15813
rect 15842 15802 15848 15804
rect 15904 15802 15928 15804
rect 15984 15802 16008 15804
rect 16064 15802 16088 15804
rect 16144 15802 16150 15804
rect 15904 15750 15906 15802
rect 16086 15750 16088 15802
rect 15842 15748 15848 15750
rect 15904 15748 15928 15750
rect 15984 15748 16008 15750
rect 16064 15748 16088 15750
rect 16144 15748 16150 15750
rect 15842 15739 16150 15748
rect 16224 15586 16252 17682
rect 16502 17436 16810 17445
rect 16502 17434 16508 17436
rect 16564 17434 16588 17436
rect 16644 17434 16668 17436
rect 16724 17434 16748 17436
rect 16804 17434 16810 17436
rect 16564 17382 16566 17434
rect 16746 17382 16748 17434
rect 16502 17380 16508 17382
rect 16564 17380 16588 17382
rect 16644 17380 16668 17382
rect 16724 17380 16748 17382
rect 16804 17380 16810 17382
rect 16502 17371 16810 17380
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 16502 16348 16810 16357
rect 16502 16346 16508 16348
rect 16564 16346 16588 16348
rect 16644 16346 16668 16348
rect 16724 16346 16748 16348
rect 16804 16346 16810 16348
rect 16564 16294 16566 16346
rect 16746 16294 16748 16346
rect 16502 16292 16508 16294
rect 16564 16292 16588 16294
rect 16644 16292 16668 16294
rect 16724 16292 16748 16294
rect 16804 16292 16810 16294
rect 16502 16283 16810 16292
rect 17052 16250 17080 16390
rect 17040 16244 17092 16250
rect 17040 16186 17092 16192
rect 16488 16040 16540 16046
rect 16488 15982 16540 15988
rect 16132 15558 16252 15586
rect 16132 15502 16160 15558
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 16120 15496 16172 15502
rect 16120 15438 16172 15444
rect 15856 15366 15884 15438
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15660 14952 15712 14958
rect 15660 14894 15712 14900
rect 15856 14890 15884 15302
rect 16132 15026 16160 15438
rect 16304 15428 16356 15434
rect 16304 15370 16356 15376
rect 16316 15162 16344 15370
rect 16500 15366 16528 15982
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17696 15745 17724 15846
rect 17682 15736 17738 15745
rect 17682 15671 17738 15680
rect 17500 15496 17552 15502
rect 17500 15438 17552 15444
rect 16488 15360 16540 15366
rect 16488 15302 16540 15308
rect 16502 15260 16810 15269
rect 16502 15258 16508 15260
rect 16564 15258 16588 15260
rect 16644 15258 16668 15260
rect 16724 15258 16748 15260
rect 16804 15258 16810 15260
rect 16564 15206 16566 15258
rect 16746 15206 16748 15258
rect 16502 15204 16508 15206
rect 16564 15204 16588 15206
rect 16644 15204 16668 15206
rect 16724 15204 16748 15206
rect 16804 15204 16810 15206
rect 16502 15195 16810 15204
rect 16304 15156 16356 15162
rect 16304 15098 16356 15104
rect 16120 15020 16172 15026
rect 16120 14962 16172 14968
rect 16396 14952 16448 14958
rect 16396 14894 16448 14900
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15660 14816 15712 14822
rect 15660 14758 15712 14764
rect 15672 14346 15700 14758
rect 15842 14716 16150 14725
rect 15842 14714 15848 14716
rect 15904 14714 15928 14716
rect 15984 14714 16008 14716
rect 16064 14714 16088 14716
rect 16144 14714 16150 14716
rect 15904 14662 15906 14714
rect 16086 14662 16088 14714
rect 15842 14660 15848 14662
rect 15904 14660 15928 14662
rect 15984 14660 16008 14662
rect 16064 14660 16088 14662
rect 16144 14660 16150 14662
rect 15842 14651 16150 14660
rect 16408 14550 16436 14894
rect 16856 14816 16908 14822
rect 16856 14758 16908 14764
rect 16396 14544 16448 14550
rect 16396 14486 16448 14492
rect 15752 14476 15804 14482
rect 15752 14418 15804 14424
rect 15660 14340 15712 14346
rect 15660 14282 15712 14288
rect 15660 13864 15712 13870
rect 15660 13806 15712 13812
rect 15568 13524 15620 13530
rect 15568 13466 15620 13472
rect 15476 13320 15528 13326
rect 15476 13262 15528 13268
rect 15488 13002 15516 13262
rect 15580 13258 15608 13466
rect 15568 13252 15620 13258
rect 15568 13194 15620 13200
rect 15672 13190 15700 13806
rect 15660 13184 15712 13190
rect 15660 13126 15712 13132
rect 15488 12974 15700 13002
rect 15200 12912 15252 12918
rect 15200 12854 15252 12860
rect 15108 12300 15160 12306
rect 15108 12242 15160 12248
rect 15200 12300 15252 12306
rect 15200 12242 15252 12248
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14924 12232 14976 12238
rect 14924 12174 14976 12180
rect 14648 11756 14700 11762
rect 14648 11698 14700 11704
rect 14844 11642 14872 12174
rect 14936 11830 14964 12174
rect 14924 11824 14976 11830
rect 14924 11766 14976 11772
rect 15016 11756 15068 11762
rect 15016 11698 15068 11704
rect 14844 11614 14964 11642
rect 14936 11286 14964 11614
rect 14924 11280 14976 11286
rect 14924 11222 14976 11228
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 14832 10668 14884 10674
rect 14832 10610 14884 10616
rect 14464 10532 14516 10538
rect 14464 10474 14516 10480
rect 14476 9926 14504 10474
rect 14556 10464 14608 10470
rect 14556 10406 14608 10412
rect 14464 9920 14516 9926
rect 14464 9862 14516 9868
rect 14568 9654 14596 10406
rect 14844 10266 14872 10610
rect 14832 10260 14884 10266
rect 14832 10202 14884 10208
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14372 8968 14424 8974
rect 14372 8910 14424 8916
rect 14280 8628 14332 8634
rect 14280 8570 14332 8576
rect 14568 8498 14596 9114
rect 14740 8968 14792 8974
rect 14740 8910 14792 8916
rect 14752 8634 14780 8910
rect 14832 8900 14884 8906
rect 14832 8842 14884 8848
rect 14740 8628 14792 8634
rect 14740 8570 14792 8576
rect 14372 8492 14424 8498
rect 14372 8434 14424 8440
rect 14556 8492 14608 8498
rect 14556 8434 14608 8440
rect 14384 8362 14412 8434
rect 14372 8356 14424 8362
rect 14372 8298 14424 8304
rect 14370 7984 14426 7993
rect 14568 7954 14596 8434
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14370 7919 14426 7928
rect 14556 7948 14608 7954
rect 14384 7886 14412 7919
rect 14556 7890 14608 7896
rect 14004 7880 14056 7886
rect 14004 7822 14056 7828
rect 14372 7880 14424 7886
rect 14372 7822 14424 7828
rect 14554 7848 14610 7857
rect 13832 7670 13952 7698
rect 13832 7562 13860 7670
rect 13544 7540 13596 7546
rect 13544 7482 13596 7488
rect 13648 7534 13860 7562
rect 13648 7410 13676 7534
rect 13912 7472 13964 7478
rect 13740 7420 13912 7426
rect 13740 7414 13964 7420
rect 13636 7404 13688 7410
rect 13636 7346 13688 7352
rect 13740 7398 13952 7414
rect 14016 7410 14044 7822
rect 14004 7404 14056 7410
rect 13636 7200 13688 7206
rect 13636 7142 13688 7148
rect 13452 6724 13504 6730
rect 13452 6666 13504 6672
rect 13268 6384 13320 6390
rect 13268 6326 13320 6332
rect 13280 5778 13308 6326
rect 13452 5840 13504 5846
rect 13452 5782 13504 5788
rect 13268 5772 13320 5778
rect 13268 5714 13320 5720
rect 13280 5370 13308 5714
rect 13360 5568 13412 5574
rect 13360 5510 13412 5516
rect 13268 5364 13320 5370
rect 13268 5306 13320 5312
rect 13176 5228 13228 5234
rect 13176 5170 13228 5176
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 13096 4078 13124 5102
rect 13084 4072 13136 4078
rect 13084 4014 13136 4020
rect 13096 3482 13124 4014
rect 13096 3466 13216 3482
rect 13096 3460 13228 3466
rect 13096 3454 13176 3460
rect 13176 3402 13228 3408
rect 13372 3346 13400 5510
rect 13464 4622 13492 5782
rect 13544 5772 13596 5778
rect 13544 5714 13596 5720
rect 13556 5642 13584 5714
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13544 5024 13596 5030
rect 13544 4966 13596 4972
rect 13556 4826 13584 4966
rect 13544 4820 13596 4826
rect 13544 4762 13596 4768
rect 13648 4622 13676 7142
rect 13740 6662 13768 7398
rect 14004 7346 14056 7352
rect 13728 6656 13780 6662
rect 13728 6598 13780 6604
rect 14016 6361 14044 7346
rect 14280 7336 14332 7342
rect 14280 7278 14332 7284
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14096 6860 14148 6866
rect 14096 6802 14148 6808
rect 14002 6352 14058 6361
rect 14002 6287 14058 6296
rect 14108 6254 14136 6802
rect 14096 6248 14148 6254
rect 14096 6190 14148 6196
rect 13728 5228 13780 5234
rect 13728 5170 13780 5176
rect 13820 5228 13872 5234
rect 13820 5170 13872 5176
rect 13452 4616 13504 4622
rect 13452 4558 13504 4564
rect 13636 4616 13688 4622
rect 13636 4558 13688 4564
rect 13452 4480 13504 4486
rect 13452 4422 13504 4428
rect 13464 4078 13492 4422
rect 13544 4276 13596 4282
rect 13544 4218 13596 4224
rect 13452 4072 13504 4078
rect 13452 4014 13504 4020
rect 13556 3534 13584 4218
rect 13740 4146 13768 5170
rect 13832 4690 13860 5170
rect 14200 4690 14228 7142
rect 14292 6730 14320 7278
rect 14384 6798 14412 7822
rect 14554 7783 14610 7792
rect 14464 7540 14516 7546
rect 14464 7482 14516 7488
rect 14476 6798 14504 7482
rect 14568 7342 14596 7783
rect 14648 7744 14700 7750
rect 14648 7686 14700 7692
rect 14660 7342 14688 7686
rect 14556 7336 14608 7342
rect 14556 7278 14608 7284
rect 14648 7336 14700 7342
rect 14648 7278 14700 7284
rect 14372 6792 14424 6798
rect 14372 6734 14424 6740
rect 14464 6792 14516 6798
rect 14464 6734 14516 6740
rect 14280 6724 14332 6730
rect 14280 6666 14332 6672
rect 14370 5808 14426 5817
rect 14370 5743 14372 5752
rect 14424 5743 14426 5752
rect 14372 5714 14424 5720
rect 13820 4684 13872 4690
rect 13820 4626 13872 4632
rect 14188 4684 14240 4690
rect 14188 4626 14240 4632
rect 13832 4146 13860 4626
rect 14004 4548 14056 4554
rect 14004 4490 14056 4496
rect 14016 4146 14044 4490
rect 14384 4486 14412 5714
rect 14568 5710 14596 7278
rect 14660 6916 14688 7278
rect 14752 7206 14780 8366
rect 14740 7200 14792 7206
rect 14740 7142 14792 7148
rect 14844 7002 14872 8842
rect 14936 8362 14964 11222
rect 15028 11218 15056 11698
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 15028 10033 15056 11154
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 10538 15148 10950
rect 15108 10532 15160 10538
rect 15108 10474 15160 10480
rect 15212 10130 15240 12242
rect 15672 12170 15700 12974
rect 15660 12164 15712 12170
rect 15660 12106 15712 12112
rect 15764 11830 15792 14418
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 15842 13628 16150 13637
rect 15842 13626 15848 13628
rect 15904 13626 15928 13628
rect 15984 13626 16008 13628
rect 16064 13626 16088 13628
rect 16144 13626 16150 13628
rect 15904 13574 15906 13626
rect 16086 13574 16088 13626
rect 15842 13572 15848 13574
rect 15904 13572 15928 13574
rect 15984 13572 16008 13574
rect 16064 13572 16088 13574
rect 16144 13572 16150 13574
rect 15842 13563 16150 13572
rect 16224 13530 16252 14214
rect 16408 14074 16436 14486
rect 16868 14346 16896 14758
rect 16946 14376 17002 14385
rect 16856 14340 16908 14346
rect 16946 14311 17002 14320
rect 16856 14282 16908 14288
rect 16502 14172 16810 14181
rect 16502 14170 16508 14172
rect 16564 14170 16588 14172
rect 16644 14170 16668 14172
rect 16724 14170 16748 14172
rect 16804 14170 16810 14172
rect 16564 14118 16566 14170
rect 16746 14118 16748 14170
rect 16502 14116 16508 14118
rect 16564 14116 16588 14118
rect 16644 14116 16668 14118
rect 16724 14116 16748 14118
rect 16804 14116 16810 14118
rect 16502 14107 16810 14116
rect 16960 14074 16988 14311
rect 16396 14068 16448 14074
rect 16396 14010 16448 14016
rect 16948 14068 17000 14074
rect 16948 14010 17000 14016
rect 16304 14000 16356 14006
rect 16304 13942 16356 13948
rect 16212 13524 16264 13530
rect 16212 13466 16264 13472
rect 15842 12540 16150 12549
rect 15842 12538 15848 12540
rect 15904 12538 15928 12540
rect 15984 12538 16008 12540
rect 16064 12538 16088 12540
rect 16144 12538 16150 12540
rect 15904 12486 15906 12538
rect 16086 12486 16088 12538
rect 15842 12484 15848 12486
rect 15904 12484 15928 12486
rect 15984 12484 16008 12486
rect 16064 12484 16088 12486
rect 16144 12484 16150 12486
rect 15842 12475 16150 12484
rect 16224 12322 16252 13466
rect 16316 12594 16344 13942
rect 17132 13728 17184 13734
rect 17132 13670 17184 13676
rect 17144 13326 17172 13670
rect 17512 13462 17540 15438
rect 17684 15360 17736 15366
rect 17684 15302 17736 15308
rect 17696 15065 17724 15302
rect 17682 15056 17738 15065
rect 17682 14991 17738 15000
rect 17776 15020 17828 15026
rect 17776 14962 17828 14968
rect 17592 14816 17644 14822
rect 17592 14758 17644 14764
rect 17604 14346 17632 14758
rect 17788 14618 17816 14962
rect 17776 14612 17828 14618
rect 17776 14554 17828 14560
rect 17592 14340 17644 14346
rect 17592 14282 17644 14288
rect 17500 13456 17552 13462
rect 17500 13398 17552 13404
rect 17224 13388 17276 13394
rect 17224 13330 17276 13336
rect 17132 13320 17184 13326
rect 17132 13262 17184 13268
rect 16502 13084 16810 13093
rect 16502 13082 16508 13084
rect 16564 13082 16588 13084
rect 16644 13082 16668 13084
rect 16724 13082 16748 13084
rect 16804 13082 16810 13084
rect 16564 13030 16566 13082
rect 16746 13030 16748 13082
rect 16502 13028 16508 13030
rect 16564 13028 16588 13030
rect 16644 13028 16668 13030
rect 16724 13028 16748 13030
rect 16804 13028 16810 13030
rect 16502 13019 16810 13028
rect 16580 12844 16632 12850
rect 16580 12786 16632 12792
rect 16488 12776 16540 12782
rect 16488 12718 16540 12724
rect 16316 12566 16436 12594
rect 16302 12472 16358 12481
rect 16408 12442 16436 12566
rect 16302 12407 16304 12416
rect 16356 12407 16358 12416
rect 16396 12436 16448 12442
rect 16304 12378 16356 12384
rect 16396 12378 16448 12384
rect 16500 12322 16528 12718
rect 16592 12481 16620 12786
rect 16672 12640 16724 12646
rect 16672 12582 16724 12588
rect 16578 12472 16634 12481
rect 16578 12407 16634 12416
rect 16224 12294 16528 12322
rect 16684 12306 16712 12582
rect 17236 12434 17264 13330
rect 17684 13252 17736 13258
rect 17684 13194 17736 13200
rect 17500 13184 17552 13190
rect 17500 13126 17552 13132
rect 17236 12406 17356 12434
rect 16672 12300 16724 12306
rect 16408 12238 16436 12294
rect 16672 12242 16724 12248
rect 16396 12232 16448 12238
rect 16396 12174 16448 12180
rect 15752 11824 15804 11830
rect 15752 11766 15804 11772
rect 16212 11688 16264 11694
rect 16212 11630 16264 11636
rect 15752 11552 15804 11558
rect 15752 11494 15804 11500
rect 15764 11082 15792 11494
rect 15842 11452 16150 11461
rect 15842 11450 15848 11452
rect 15904 11450 15928 11452
rect 15984 11450 16008 11452
rect 16064 11450 16088 11452
rect 16144 11450 16150 11452
rect 15904 11398 15906 11450
rect 16086 11398 16088 11450
rect 15842 11396 15848 11398
rect 15904 11396 15928 11398
rect 15984 11396 16008 11398
rect 16064 11396 16088 11398
rect 16144 11396 16150 11398
rect 15842 11387 16150 11396
rect 16224 11286 16252 11630
rect 16212 11280 16264 11286
rect 16212 11222 16264 11228
rect 16408 11150 16436 12174
rect 16502 11996 16810 12005
rect 16502 11994 16508 11996
rect 16564 11994 16588 11996
rect 16644 11994 16668 11996
rect 16724 11994 16748 11996
rect 16804 11994 16810 11996
rect 16564 11942 16566 11994
rect 16746 11942 16748 11994
rect 16502 11940 16508 11942
rect 16564 11940 16588 11942
rect 16644 11940 16668 11942
rect 16724 11940 16748 11942
rect 16804 11940 16810 11942
rect 16502 11931 16810 11940
rect 17132 11688 17184 11694
rect 17132 11630 17184 11636
rect 17224 11688 17276 11694
rect 17224 11630 17276 11636
rect 16396 11144 16448 11150
rect 16396 11086 16448 11092
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15568 11008 15620 11014
rect 15568 10950 15620 10956
rect 15580 10810 15608 10950
rect 15568 10804 15620 10810
rect 15568 10746 15620 10752
rect 16408 10674 16436 11086
rect 16856 11008 16908 11014
rect 16856 10950 16908 10956
rect 16502 10908 16810 10917
rect 16502 10906 16508 10908
rect 16564 10906 16588 10908
rect 16644 10906 16668 10908
rect 16724 10906 16748 10908
rect 16804 10906 16810 10908
rect 16564 10854 16566 10906
rect 16746 10854 16748 10906
rect 16502 10852 16508 10854
rect 16564 10852 16588 10854
rect 16644 10852 16668 10854
rect 16724 10852 16748 10854
rect 16804 10852 16810 10854
rect 16502 10843 16810 10852
rect 16212 10668 16264 10674
rect 16212 10610 16264 10616
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 15842 10364 16150 10373
rect 15842 10362 15848 10364
rect 15904 10362 15928 10364
rect 15984 10362 16008 10364
rect 16064 10362 16088 10364
rect 16144 10362 16150 10364
rect 15904 10310 15906 10362
rect 16086 10310 16088 10362
rect 15842 10308 15848 10310
rect 15904 10308 15928 10310
rect 15984 10308 16008 10310
rect 16064 10308 16088 10310
rect 16144 10308 16150 10310
rect 15842 10299 16150 10308
rect 16224 10266 16252 10610
rect 16672 10464 16724 10470
rect 16672 10406 16724 10412
rect 16212 10260 16264 10266
rect 16212 10202 16264 10208
rect 15200 10124 15252 10130
rect 15200 10066 15252 10072
rect 15014 10024 15070 10033
rect 15014 9959 15070 9968
rect 15016 9512 15068 9518
rect 15016 9454 15068 9460
rect 15028 8974 15056 9454
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14924 8356 14976 8362
rect 14924 8298 14976 8304
rect 14936 7449 14964 8298
rect 15028 7750 15056 8910
rect 15212 8430 15240 10066
rect 16684 10062 16712 10406
rect 16868 10130 16896 10950
rect 17144 10606 17172 11630
rect 17132 10600 17184 10606
rect 17132 10542 17184 10548
rect 16856 10124 16908 10130
rect 16856 10066 16908 10072
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16502 9820 16810 9829
rect 16502 9818 16508 9820
rect 16564 9818 16588 9820
rect 16644 9818 16668 9820
rect 16724 9818 16748 9820
rect 16804 9818 16810 9820
rect 16564 9766 16566 9818
rect 16746 9766 16748 9818
rect 16502 9764 16508 9766
rect 16564 9764 16588 9766
rect 16644 9764 16668 9766
rect 16724 9764 16748 9766
rect 16804 9764 16810 9766
rect 16502 9755 16810 9764
rect 15384 9580 15436 9586
rect 15384 9522 15436 9528
rect 15396 8906 15424 9522
rect 16304 9512 16356 9518
rect 16304 9454 16356 9460
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 15660 9444 15712 9450
rect 15660 9386 15712 9392
rect 15384 8900 15436 8906
rect 15384 8842 15436 8848
rect 15200 8424 15252 8430
rect 15200 8366 15252 8372
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 14922 7440 14978 7449
rect 14922 7375 14978 7384
rect 15108 7404 15160 7410
rect 14832 6996 14884 7002
rect 14832 6938 14884 6944
rect 14740 6928 14792 6934
rect 14660 6888 14740 6916
rect 14556 5704 14608 5710
rect 14462 5672 14518 5681
rect 14556 5646 14608 5652
rect 14462 5607 14518 5616
rect 14476 4622 14504 5607
rect 14660 5166 14688 6888
rect 14844 6905 14872 6938
rect 14740 6870 14792 6876
rect 14830 6896 14886 6905
rect 14830 6831 14886 6840
rect 14936 5914 14964 7375
rect 15108 7346 15160 7352
rect 15016 7268 15068 7274
rect 15016 7210 15068 7216
rect 15028 6322 15056 7210
rect 15016 6316 15068 6322
rect 15016 6258 15068 6264
rect 14924 5908 14976 5914
rect 14924 5850 14976 5856
rect 14832 5228 14884 5234
rect 14832 5170 14884 5176
rect 14648 5160 14700 5166
rect 14648 5102 14700 5108
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 14556 4616 14608 4622
rect 14556 4558 14608 4564
rect 14372 4480 14424 4486
rect 14372 4422 14424 4428
rect 14568 4282 14596 4558
rect 14660 4554 14688 5102
rect 14844 4826 14872 5170
rect 15120 5114 15148 7346
rect 15292 6384 15344 6390
rect 15292 6326 15344 6332
rect 15200 5568 15252 5574
rect 15200 5510 15252 5516
rect 15212 5302 15240 5510
rect 15200 5296 15252 5302
rect 15200 5238 15252 5244
rect 15120 5086 15240 5114
rect 14832 4820 14884 4826
rect 14832 4762 14884 4768
rect 14648 4548 14700 4554
rect 14648 4490 14700 4496
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 13728 4140 13780 4146
rect 13728 4082 13780 4088
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 14004 4140 14056 4146
rect 14004 4082 14056 4088
rect 13740 3602 13768 4082
rect 13728 3596 13780 3602
rect 13648 3556 13728 3584
rect 13544 3528 13596 3534
rect 13544 3470 13596 3476
rect 12820 3012 13032 3040
rect 13096 3318 13400 3346
rect 12072 2508 12124 2514
rect 12072 2450 12124 2456
rect 12716 2440 12768 2446
rect 12820 2428 12848 3012
rect 13096 2938 13124 3318
rect 13176 3188 13228 3194
rect 13176 3130 13228 3136
rect 12912 2910 13124 2938
rect 12912 2446 12940 2910
rect 13188 2446 13216 3130
rect 13556 2582 13584 3470
rect 13648 2854 13676 3556
rect 13728 3538 13780 3544
rect 14096 3528 14148 3534
rect 14096 3470 14148 3476
rect 13636 2848 13688 2854
rect 13636 2790 13688 2796
rect 14108 2650 14136 3470
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 14292 3058 14320 3334
rect 14660 3058 14688 4490
rect 15212 4146 15240 5086
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15304 3942 15332 6326
rect 15396 5846 15424 8842
rect 15568 8832 15620 8838
rect 15568 8774 15620 8780
rect 15580 8498 15608 8774
rect 15672 8634 15700 9386
rect 15842 9276 16150 9285
rect 15842 9274 15848 9276
rect 15904 9274 15928 9276
rect 15984 9274 16008 9276
rect 16064 9274 16088 9276
rect 16144 9274 16150 9276
rect 15904 9222 15906 9274
rect 16086 9222 16088 9274
rect 15842 9220 15848 9222
rect 15904 9220 15928 9222
rect 15984 9220 16008 9222
rect 16064 9220 16088 9222
rect 16144 9220 16150 9222
rect 15842 9211 16150 9220
rect 15752 8900 15804 8906
rect 15752 8842 15804 8848
rect 15764 8634 15792 8842
rect 15660 8628 15712 8634
rect 15660 8570 15712 8576
rect 15752 8628 15804 8634
rect 15752 8570 15804 8576
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15476 8424 15528 8430
rect 15476 8366 15528 8372
rect 15488 6866 15516 8366
rect 15476 6860 15528 6866
rect 15476 6802 15528 6808
rect 15580 6390 15608 8434
rect 15764 6916 15792 8570
rect 16212 8492 16264 8498
rect 16212 8434 16264 8440
rect 15842 8188 16150 8197
rect 15842 8186 15848 8188
rect 15904 8186 15928 8188
rect 15984 8186 16008 8188
rect 16064 8186 16088 8188
rect 16144 8186 16150 8188
rect 15904 8134 15906 8186
rect 16086 8134 16088 8186
rect 15842 8132 15848 8134
rect 15904 8132 15928 8134
rect 15984 8132 16008 8134
rect 16064 8132 16088 8134
rect 16144 8132 16150 8134
rect 15842 8123 16150 8132
rect 15842 7100 16150 7109
rect 15842 7098 15848 7100
rect 15904 7098 15928 7100
rect 15984 7098 16008 7100
rect 16064 7098 16088 7100
rect 16144 7098 16150 7100
rect 15904 7046 15906 7098
rect 16086 7046 16088 7098
rect 15842 7044 15848 7046
rect 15904 7044 15928 7046
rect 15984 7044 16008 7046
rect 16064 7044 16088 7046
rect 16144 7044 16150 7046
rect 15842 7035 16150 7044
rect 15764 6888 15884 6916
rect 15660 6656 15712 6662
rect 15660 6598 15712 6604
rect 15752 6656 15804 6662
rect 15752 6598 15804 6604
rect 15672 6458 15700 6598
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15568 6384 15620 6390
rect 15568 6326 15620 6332
rect 15476 6248 15528 6254
rect 15476 6190 15528 6196
rect 15384 5840 15436 5846
rect 15384 5782 15436 5788
rect 15384 5704 15436 5710
rect 15384 5646 15436 5652
rect 15396 4826 15424 5646
rect 15384 4820 15436 4826
rect 15384 4762 15436 4768
rect 15488 4570 15516 6190
rect 15764 5930 15792 6598
rect 15856 6254 15884 6888
rect 16224 6662 16252 8434
rect 16316 8090 16344 9454
rect 16408 9178 16436 9454
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16396 9172 16448 9178
rect 16396 9114 16448 9120
rect 16500 8974 16528 9318
rect 17236 9042 17264 11630
rect 17328 10606 17356 12406
rect 17512 11762 17540 13126
rect 17696 13025 17724 13194
rect 17682 13016 17738 13025
rect 17682 12951 17738 12960
rect 17684 12164 17736 12170
rect 17684 12106 17736 12112
rect 17696 11898 17724 12106
rect 17684 11892 17736 11898
rect 17684 11834 17736 11840
rect 17500 11756 17552 11762
rect 17500 11698 17552 11704
rect 17500 10668 17552 10674
rect 17500 10610 17552 10616
rect 17684 10668 17736 10674
rect 17684 10610 17736 10616
rect 17316 10600 17368 10606
rect 17316 10542 17368 10548
rect 17224 9036 17276 9042
rect 17224 8978 17276 8984
rect 16488 8968 16540 8974
rect 16488 8910 16540 8916
rect 16502 8732 16810 8741
rect 16502 8730 16508 8732
rect 16564 8730 16588 8732
rect 16644 8730 16668 8732
rect 16724 8730 16748 8732
rect 16804 8730 16810 8732
rect 16564 8678 16566 8730
rect 16746 8678 16748 8730
rect 16502 8676 16508 8678
rect 16564 8676 16588 8678
rect 16644 8676 16668 8678
rect 16724 8676 16748 8678
rect 16804 8676 16810 8678
rect 16502 8667 16810 8676
rect 17328 8634 17356 10542
rect 17512 10266 17540 10610
rect 17696 10305 17724 10610
rect 17682 10296 17738 10305
rect 17500 10260 17552 10266
rect 17682 10231 17738 10240
rect 17500 10202 17552 10208
rect 17500 8832 17552 8838
rect 17500 8774 17552 8780
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 16948 8424 17000 8430
rect 16948 8366 17000 8372
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16304 8084 16356 8090
rect 16304 8026 16356 8032
rect 16316 7546 16344 8026
rect 16304 7540 16356 7546
rect 16304 7482 16356 7488
rect 16408 7410 16436 8298
rect 16960 8265 16988 8366
rect 16946 8256 17002 8265
rect 16946 8191 17002 8200
rect 17512 7818 17540 8774
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 16502 7644 16810 7653
rect 16502 7642 16508 7644
rect 16564 7642 16588 7644
rect 16644 7642 16668 7644
rect 16724 7642 16748 7644
rect 16804 7642 16810 7644
rect 16564 7590 16566 7642
rect 16746 7590 16748 7642
rect 16502 7588 16508 7590
rect 16564 7588 16588 7590
rect 16644 7588 16668 7590
rect 16724 7588 16748 7590
rect 16804 7588 16810 7590
rect 16502 7579 16810 7588
rect 17774 7576 17830 7585
rect 17774 7511 17830 7520
rect 17788 7410 17816 7511
rect 16396 7404 16448 7410
rect 16396 7346 16448 7352
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17774 6896 17830 6905
rect 17774 6831 17830 6840
rect 16396 6724 16448 6730
rect 16396 6666 16448 6672
rect 16856 6724 16908 6730
rect 16856 6666 16908 6672
rect 16212 6656 16264 6662
rect 16212 6598 16264 6604
rect 16304 6316 16356 6322
rect 16304 6258 16356 6264
rect 15844 6248 15896 6254
rect 15844 6190 15896 6196
rect 15842 6012 16150 6021
rect 15842 6010 15848 6012
rect 15904 6010 15928 6012
rect 15984 6010 16008 6012
rect 16064 6010 16088 6012
rect 16144 6010 16150 6012
rect 15904 5958 15906 6010
rect 16086 5958 16088 6010
rect 15842 5956 15848 5958
rect 15904 5956 15928 5958
rect 15984 5956 16008 5958
rect 16064 5956 16088 5958
rect 16144 5956 16150 5958
rect 15842 5947 16150 5956
rect 15396 4542 15516 4570
rect 15580 5902 15792 5930
rect 15396 4282 15424 4542
rect 15580 4486 15608 5902
rect 15764 5794 15792 5902
rect 15764 5778 15884 5794
rect 15660 5772 15712 5778
rect 15764 5772 15896 5778
rect 15764 5766 15844 5772
rect 15660 5714 15712 5720
rect 15844 5714 15896 5720
rect 15672 4486 15700 5714
rect 15752 5636 15804 5642
rect 15752 5578 15804 5584
rect 15568 4480 15620 4486
rect 15488 4428 15568 4434
rect 15488 4422 15620 4428
rect 15660 4480 15712 4486
rect 15660 4422 15712 4428
rect 15488 4406 15608 4422
rect 15384 4276 15436 4282
rect 15384 4218 15436 4224
rect 15488 4214 15516 4406
rect 15476 4208 15528 4214
rect 15476 4150 15528 4156
rect 15672 4078 15700 4422
rect 15764 4146 15792 5578
rect 16212 5024 16264 5030
rect 16212 4966 16264 4972
rect 15842 4924 16150 4933
rect 15842 4922 15848 4924
rect 15904 4922 15928 4924
rect 15984 4922 16008 4924
rect 16064 4922 16088 4924
rect 16144 4922 16150 4924
rect 15904 4870 15906 4922
rect 16086 4870 16088 4922
rect 15842 4868 15848 4870
rect 15904 4868 15928 4870
rect 15984 4868 16008 4870
rect 16064 4868 16088 4870
rect 16144 4868 16150 4870
rect 15842 4859 16150 4868
rect 16224 4758 16252 4966
rect 16212 4752 16264 4758
rect 16212 4694 16264 4700
rect 15844 4684 15896 4690
rect 15844 4626 15896 4632
rect 15856 4282 15884 4626
rect 15844 4276 15896 4282
rect 15844 4218 15896 4224
rect 16316 4146 16344 6258
rect 16408 6254 16436 6666
rect 16502 6556 16810 6565
rect 16502 6554 16508 6556
rect 16564 6554 16588 6556
rect 16644 6554 16668 6556
rect 16724 6554 16748 6556
rect 16804 6554 16810 6556
rect 16564 6502 16566 6554
rect 16746 6502 16748 6554
rect 16502 6500 16508 6502
rect 16564 6500 16588 6502
rect 16644 6500 16668 6502
rect 16724 6500 16748 6502
rect 16804 6500 16810 6502
rect 16502 6491 16810 6500
rect 16868 6458 16896 6666
rect 17500 6656 17552 6662
rect 17500 6598 17552 6604
rect 16856 6452 16908 6458
rect 16856 6394 16908 6400
rect 16396 6248 16448 6254
rect 16396 6190 16448 6196
rect 16408 4214 16436 6190
rect 17040 5568 17092 5574
rect 17040 5510 17092 5516
rect 16502 5468 16810 5477
rect 16502 5466 16508 5468
rect 16564 5466 16588 5468
rect 16644 5466 16668 5468
rect 16724 5466 16748 5468
rect 16804 5466 16810 5468
rect 16564 5414 16566 5466
rect 16746 5414 16748 5466
rect 16502 5412 16508 5414
rect 16564 5412 16588 5414
rect 16644 5412 16668 5414
rect 16724 5412 16748 5414
rect 16804 5412 16810 5414
rect 16502 5403 16810 5412
rect 17052 4554 17080 5510
rect 17040 4548 17092 4554
rect 17040 4490 17092 4496
rect 16502 4380 16810 4389
rect 16502 4378 16508 4380
rect 16564 4378 16588 4380
rect 16644 4378 16668 4380
rect 16724 4378 16748 4380
rect 16804 4378 16810 4380
rect 16564 4326 16566 4378
rect 16746 4326 16748 4378
rect 16502 4324 16508 4326
rect 16564 4324 16588 4326
rect 16644 4324 16668 4326
rect 16724 4324 16748 4326
rect 16804 4324 16810 4326
rect 16502 4315 16810 4324
rect 16396 4208 16448 4214
rect 16396 4150 16448 4156
rect 17512 4146 17540 6598
rect 17788 6322 17816 6831
rect 17776 6316 17828 6322
rect 17776 6258 17828 6264
rect 17774 6216 17830 6225
rect 17774 6151 17830 6160
rect 17788 5778 17816 6151
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17682 5536 17738 5545
rect 17682 5471 17738 5480
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 17604 4865 17632 4966
rect 17590 4856 17646 4865
rect 17696 4826 17724 5471
rect 17590 4791 17646 4800
rect 17684 4820 17736 4826
rect 17684 4762 17736 4768
rect 15752 4140 15804 4146
rect 15752 4082 15804 4088
rect 16304 4140 16356 4146
rect 16304 4082 16356 4088
rect 17500 4140 17552 4146
rect 17500 4082 17552 4088
rect 15660 4072 15712 4078
rect 15660 4014 15712 4020
rect 15292 3936 15344 3942
rect 15292 3878 15344 3884
rect 15304 3602 15332 3878
rect 15842 3836 16150 3845
rect 15842 3834 15848 3836
rect 15904 3834 15928 3836
rect 15984 3834 16008 3836
rect 16064 3834 16088 3836
rect 16144 3834 16150 3836
rect 15904 3782 15906 3834
rect 16086 3782 16088 3834
rect 15842 3780 15848 3782
rect 15904 3780 15928 3782
rect 15984 3780 16008 3782
rect 16064 3780 16088 3782
rect 16144 3780 16150 3782
rect 15842 3771 16150 3780
rect 15292 3596 15344 3602
rect 15292 3538 15344 3544
rect 15304 3398 15332 3538
rect 16028 3528 16080 3534
rect 16028 3470 16080 3476
rect 17682 3496 17738 3505
rect 14740 3392 14792 3398
rect 14740 3334 14792 3340
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 15292 3392 15344 3398
rect 15292 3334 15344 3340
rect 14752 3126 14780 3334
rect 14740 3120 14792 3126
rect 14740 3062 14792 3068
rect 14280 3052 14332 3058
rect 14280 2994 14332 3000
rect 14648 3052 14700 3058
rect 14648 2994 14700 3000
rect 14646 2952 14702 2961
rect 14646 2887 14702 2896
rect 14096 2644 14148 2650
rect 14096 2586 14148 2592
rect 13544 2576 13596 2582
rect 13544 2518 13596 2524
rect 14660 2514 14688 2887
rect 14936 2582 14964 3334
rect 16040 3194 16068 3470
rect 17682 3431 17684 3440
rect 17736 3431 17738 3440
rect 17684 3402 17736 3408
rect 16502 3292 16810 3301
rect 16502 3290 16508 3292
rect 16564 3290 16588 3292
rect 16644 3290 16668 3292
rect 16724 3290 16748 3292
rect 16804 3290 16810 3292
rect 16564 3238 16566 3290
rect 16746 3238 16748 3290
rect 16502 3236 16508 3238
rect 16564 3236 16588 3238
rect 16644 3236 16668 3238
rect 16724 3236 16748 3238
rect 16804 3236 16810 3238
rect 16502 3227 16810 3236
rect 16028 3188 16080 3194
rect 16028 3130 16080 3136
rect 15842 2748 16150 2757
rect 15842 2746 15848 2748
rect 15904 2746 15928 2748
rect 15984 2746 16008 2748
rect 16064 2746 16088 2748
rect 16144 2746 16150 2748
rect 15904 2694 15906 2746
rect 16086 2694 16088 2746
rect 15842 2692 15848 2694
rect 15904 2692 15928 2694
rect 15984 2692 16008 2694
rect 16064 2692 16088 2694
rect 16144 2692 16150 2694
rect 15842 2683 16150 2692
rect 14924 2576 14976 2582
rect 14924 2518 14976 2524
rect 14648 2508 14700 2514
rect 14648 2450 14700 2456
rect 12768 2400 12848 2428
rect 12900 2440 12952 2446
rect 12716 2382 12768 2388
rect 12900 2382 12952 2388
rect 13176 2440 13228 2446
rect 13176 2382 13228 2388
rect 12164 2372 12216 2378
rect 12164 2314 12216 2320
rect 12176 1170 12204 2314
rect 12247 2204 12555 2213
rect 12247 2202 12253 2204
rect 12309 2202 12333 2204
rect 12389 2202 12413 2204
rect 12469 2202 12493 2204
rect 12549 2202 12555 2204
rect 12309 2150 12311 2202
rect 12491 2150 12493 2202
rect 12247 2148 12253 2150
rect 12309 2148 12333 2150
rect 12389 2148 12413 2150
rect 12469 2148 12493 2150
rect 12549 2148 12555 2150
rect 12247 2139 12555 2148
rect 16502 2204 16810 2213
rect 16502 2202 16508 2204
rect 16564 2202 16588 2204
rect 16644 2202 16668 2204
rect 16724 2202 16748 2204
rect 16804 2202 16810 2204
rect 16564 2150 16566 2202
rect 16746 2150 16748 2202
rect 16502 2148 16508 2150
rect 16564 2148 16588 2150
rect 16644 2148 16668 2150
rect 16724 2148 16748 2150
rect 16804 2148 16810 2150
rect 16502 2139 16810 2148
rect 12176 1142 12296 1170
rect 12268 800 12296 1142
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11610 0 11666 800
rect 12254 0 12310 800
<< via2 >>
rect 3083 19066 3139 19068
rect 3163 19066 3219 19068
rect 3243 19066 3299 19068
rect 3323 19066 3379 19068
rect 3083 19014 3129 19066
rect 3129 19014 3139 19066
rect 3163 19014 3193 19066
rect 3193 19014 3205 19066
rect 3205 19014 3219 19066
rect 3243 19014 3257 19066
rect 3257 19014 3269 19066
rect 3269 19014 3299 19066
rect 3323 19014 3333 19066
rect 3333 19014 3379 19066
rect 3083 19012 3139 19014
rect 3163 19012 3219 19014
rect 3243 19012 3299 19014
rect 3323 19012 3379 19014
rect 7338 19066 7394 19068
rect 7418 19066 7474 19068
rect 7498 19066 7554 19068
rect 7578 19066 7634 19068
rect 7338 19014 7384 19066
rect 7384 19014 7394 19066
rect 7418 19014 7448 19066
rect 7448 19014 7460 19066
rect 7460 19014 7474 19066
rect 7498 19014 7512 19066
rect 7512 19014 7524 19066
rect 7524 19014 7554 19066
rect 7578 19014 7588 19066
rect 7588 19014 7634 19066
rect 7338 19012 7394 19014
rect 7418 19012 7474 19014
rect 7498 19012 7554 19014
rect 7578 19012 7634 19014
rect 3743 18522 3799 18524
rect 3823 18522 3879 18524
rect 3903 18522 3959 18524
rect 3983 18522 4039 18524
rect 3743 18470 3789 18522
rect 3789 18470 3799 18522
rect 3823 18470 3853 18522
rect 3853 18470 3865 18522
rect 3865 18470 3879 18522
rect 3903 18470 3917 18522
rect 3917 18470 3929 18522
rect 3929 18470 3959 18522
rect 3983 18470 3993 18522
rect 3993 18470 4039 18522
rect 3743 18468 3799 18470
rect 3823 18468 3879 18470
rect 3903 18468 3959 18470
rect 3983 18468 4039 18470
rect 3083 17978 3139 17980
rect 3163 17978 3219 17980
rect 3243 17978 3299 17980
rect 3323 17978 3379 17980
rect 3083 17926 3129 17978
rect 3129 17926 3139 17978
rect 3163 17926 3193 17978
rect 3193 17926 3205 17978
rect 3205 17926 3219 17978
rect 3243 17926 3257 17978
rect 3257 17926 3269 17978
rect 3269 17926 3299 17978
rect 3323 17926 3333 17978
rect 3333 17926 3379 17978
rect 3083 17924 3139 17926
rect 3163 17924 3219 17926
rect 3243 17924 3299 17926
rect 3323 17924 3379 17926
rect 7338 17978 7394 17980
rect 7418 17978 7474 17980
rect 7498 17978 7554 17980
rect 7578 17978 7634 17980
rect 7338 17926 7384 17978
rect 7384 17926 7394 17978
rect 7418 17926 7448 17978
rect 7448 17926 7460 17978
rect 7460 17926 7474 17978
rect 7498 17926 7512 17978
rect 7512 17926 7524 17978
rect 7524 17926 7554 17978
rect 7578 17926 7588 17978
rect 7588 17926 7634 17978
rect 7338 17924 7394 17926
rect 7418 17924 7474 17926
rect 7498 17924 7554 17926
rect 7578 17924 7634 17926
rect 3743 17434 3799 17436
rect 3823 17434 3879 17436
rect 3903 17434 3959 17436
rect 3983 17434 4039 17436
rect 3743 17382 3789 17434
rect 3789 17382 3799 17434
rect 3823 17382 3853 17434
rect 3853 17382 3865 17434
rect 3865 17382 3879 17434
rect 3903 17382 3917 17434
rect 3917 17382 3929 17434
rect 3929 17382 3959 17434
rect 3983 17382 3993 17434
rect 3993 17382 4039 17434
rect 3743 17380 3799 17382
rect 3823 17380 3879 17382
rect 3903 17380 3959 17382
rect 3983 17380 4039 17382
rect 846 16516 902 16552
rect 846 16496 848 16516
rect 848 16496 900 16516
rect 900 16496 902 16516
rect 3083 16890 3139 16892
rect 3163 16890 3219 16892
rect 3243 16890 3299 16892
rect 3323 16890 3379 16892
rect 3083 16838 3129 16890
rect 3129 16838 3139 16890
rect 3163 16838 3193 16890
rect 3193 16838 3205 16890
rect 3205 16838 3219 16890
rect 3243 16838 3257 16890
rect 3257 16838 3269 16890
rect 3269 16838 3299 16890
rect 3323 16838 3333 16890
rect 3333 16838 3379 16890
rect 3083 16836 3139 16838
rect 3163 16836 3219 16838
rect 3243 16836 3299 16838
rect 3323 16836 3379 16838
rect 7998 18522 8054 18524
rect 8078 18522 8134 18524
rect 8158 18522 8214 18524
rect 8238 18522 8294 18524
rect 7998 18470 8044 18522
rect 8044 18470 8054 18522
rect 8078 18470 8108 18522
rect 8108 18470 8120 18522
rect 8120 18470 8134 18522
rect 8158 18470 8172 18522
rect 8172 18470 8184 18522
rect 8184 18470 8214 18522
rect 8238 18470 8248 18522
rect 8248 18470 8294 18522
rect 7998 18468 8054 18470
rect 8078 18468 8134 18470
rect 8158 18468 8214 18470
rect 8238 18468 8294 18470
rect 3743 16346 3799 16348
rect 3823 16346 3879 16348
rect 3903 16346 3959 16348
rect 3983 16346 4039 16348
rect 3743 16294 3789 16346
rect 3789 16294 3799 16346
rect 3823 16294 3853 16346
rect 3853 16294 3865 16346
rect 3865 16294 3879 16346
rect 3903 16294 3917 16346
rect 3917 16294 3929 16346
rect 3929 16294 3959 16346
rect 3983 16294 3993 16346
rect 3993 16294 4039 16346
rect 3743 16292 3799 16294
rect 3823 16292 3879 16294
rect 3903 16292 3959 16294
rect 3983 16292 4039 16294
rect 1490 15000 1546 15056
rect 846 14492 848 14512
rect 848 14492 900 14512
rect 900 14492 902 14512
rect 846 14456 902 14492
rect 1030 12960 1086 13016
rect 1306 12280 1362 12336
rect 3083 15802 3139 15804
rect 3163 15802 3219 15804
rect 3243 15802 3299 15804
rect 3323 15802 3379 15804
rect 3083 15750 3129 15802
rect 3129 15750 3139 15802
rect 3163 15750 3193 15802
rect 3193 15750 3205 15802
rect 3205 15750 3219 15802
rect 3243 15750 3257 15802
rect 3257 15750 3269 15802
rect 3269 15750 3299 15802
rect 3323 15750 3333 15802
rect 3333 15750 3379 15802
rect 3083 15748 3139 15750
rect 3163 15748 3219 15750
rect 3243 15748 3299 15750
rect 3323 15748 3379 15750
rect 7998 17434 8054 17436
rect 8078 17434 8134 17436
rect 8158 17434 8214 17436
rect 8238 17434 8294 17436
rect 7998 17382 8044 17434
rect 8044 17382 8054 17434
rect 8078 17382 8108 17434
rect 8108 17382 8120 17434
rect 8120 17382 8134 17434
rect 8158 17382 8172 17434
rect 8172 17382 8184 17434
rect 8184 17382 8214 17434
rect 8238 17382 8248 17434
rect 8248 17382 8294 17434
rect 7998 17380 8054 17382
rect 8078 17380 8134 17382
rect 8158 17380 8214 17382
rect 8238 17380 8294 17382
rect 3743 15258 3799 15260
rect 3823 15258 3879 15260
rect 3903 15258 3959 15260
rect 3983 15258 4039 15260
rect 3743 15206 3789 15258
rect 3789 15206 3799 15258
rect 3823 15206 3853 15258
rect 3853 15206 3865 15258
rect 3865 15206 3879 15258
rect 3903 15206 3917 15258
rect 3917 15206 3929 15258
rect 3929 15206 3959 15258
rect 3983 15206 3993 15258
rect 3993 15206 4039 15258
rect 3743 15204 3799 15206
rect 3823 15204 3879 15206
rect 3903 15204 3959 15206
rect 3983 15204 4039 15206
rect 3083 14714 3139 14716
rect 3163 14714 3219 14716
rect 3243 14714 3299 14716
rect 3323 14714 3379 14716
rect 3083 14662 3129 14714
rect 3129 14662 3139 14714
rect 3163 14662 3193 14714
rect 3193 14662 3205 14714
rect 3205 14662 3219 14714
rect 3243 14662 3257 14714
rect 3257 14662 3269 14714
rect 3269 14662 3299 14714
rect 3323 14662 3333 14714
rect 3333 14662 3379 14714
rect 3083 14660 3139 14662
rect 3163 14660 3219 14662
rect 3243 14660 3299 14662
rect 3323 14660 3379 14662
rect 1490 10920 1546 10976
rect 1214 10260 1270 10296
rect 1214 10240 1216 10260
rect 1216 10240 1268 10260
rect 1268 10240 1270 10260
rect 3083 13626 3139 13628
rect 3163 13626 3219 13628
rect 3243 13626 3299 13628
rect 3323 13626 3379 13628
rect 3083 13574 3129 13626
rect 3129 13574 3139 13626
rect 3163 13574 3193 13626
rect 3193 13574 3205 13626
rect 3205 13574 3219 13626
rect 3243 13574 3257 13626
rect 3257 13574 3269 13626
rect 3269 13574 3299 13626
rect 3323 13574 3333 13626
rect 3333 13574 3379 13626
rect 3083 13572 3139 13574
rect 3163 13572 3219 13574
rect 3243 13572 3299 13574
rect 3323 13572 3379 13574
rect 3743 14170 3799 14172
rect 3823 14170 3879 14172
rect 3903 14170 3959 14172
rect 3983 14170 4039 14172
rect 3743 14118 3789 14170
rect 3789 14118 3799 14170
rect 3823 14118 3853 14170
rect 3853 14118 3865 14170
rect 3865 14118 3879 14170
rect 3903 14118 3917 14170
rect 3917 14118 3929 14170
rect 3929 14118 3959 14170
rect 3983 14118 3993 14170
rect 3993 14118 4039 14170
rect 3743 14116 3799 14118
rect 3823 14116 3879 14118
rect 3903 14116 3959 14118
rect 3983 14116 4039 14118
rect 3743 13082 3799 13084
rect 3823 13082 3879 13084
rect 3903 13082 3959 13084
rect 3983 13082 4039 13084
rect 3743 13030 3789 13082
rect 3789 13030 3799 13082
rect 3823 13030 3853 13082
rect 3853 13030 3865 13082
rect 3865 13030 3879 13082
rect 3903 13030 3917 13082
rect 3917 13030 3929 13082
rect 3929 13030 3959 13082
rect 3983 13030 3993 13082
rect 3993 13030 4039 13082
rect 3743 13028 3799 13030
rect 3823 13028 3879 13030
rect 3903 13028 3959 13030
rect 3983 13028 4039 13030
rect 3083 12538 3139 12540
rect 3163 12538 3219 12540
rect 3243 12538 3299 12540
rect 3323 12538 3379 12540
rect 3083 12486 3129 12538
rect 3129 12486 3139 12538
rect 3163 12486 3193 12538
rect 3193 12486 3205 12538
rect 3205 12486 3219 12538
rect 3243 12486 3257 12538
rect 3257 12486 3269 12538
rect 3269 12486 3299 12538
rect 3323 12486 3333 12538
rect 3333 12486 3379 12538
rect 3083 12484 3139 12486
rect 3163 12484 3219 12486
rect 3243 12484 3299 12486
rect 3323 12484 3379 12486
rect 7338 16890 7394 16892
rect 7418 16890 7474 16892
rect 7498 16890 7554 16892
rect 7578 16890 7634 16892
rect 7338 16838 7384 16890
rect 7384 16838 7394 16890
rect 7418 16838 7448 16890
rect 7448 16838 7460 16890
rect 7460 16838 7474 16890
rect 7498 16838 7512 16890
rect 7512 16838 7524 16890
rect 7524 16838 7554 16890
rect 7578 16838 7588 16890
rect 7588 16838 7634 16890
rect 7338 16836 7394 16838
rect 7418 16836 7474 16838
rect 7498 16836 7554 16838
rect 7578 16836 7634 16838
rect 3743 11994 3799 11996
rect 3823 11994 3879 11996
rect 3903 11994 3959 11996
rect 3983 11994 4039 11996
rect 3743 11942 3789 11994
rect 3789 11942 3799 11994
rect 3823 11942 3853 11994
rect 3853 11942 3865 11994
rect 3865 11942 3879 11994
rect 3903 11942 3917 11994
rect 3917 11942 3929 11994
rect 3929 11942 3959 11994
rect 3983 11942 3993 11994
rect 3993 11942 4039 11994
rect 3743 11940 3799 11942
rect 3823 11940 3879 11942
rect 3903 11940 3959 11942
rect 3983 11940 4039 11942
rect 3083 11450 3139 11452
rect 3163 11450 3219 11452
rect 3243 11450 3299 11452
rect 3323 11450 3379 11452
rect 3083 11398 3129 11450
rect 3129 11398 3139 11450
rect 3163 11398 3193 11450
rect 3193 11398 3205 11450
rect 3205 11398 3219 11450
rect 3243 11398 3257 11450
rect 3257 11398 3269 11450
rect 3269 11398 3299 11450
rect 3323 11398 3333 11450
rect 3333 11398 3379 11450
rect 3083 11396 3139 11398
rect 3163 11396 3219 11398
rect 3243 11396 3299 11398
rect 3323 11396 3379 11398
rect 1858 9560 1914 9616
rect 3743 10906 3799 10908
rect 3823 10906 3879 10908
rect 3903 10906 3959 10908
rect 3983 10906 4039 10908
rect 3743 10854 3789 10906
rect 3789 10854 3799 10906
rect 3823 10854 3853 10906
rect 3853 10854 3865 10906
rect 3865 10854 3879 10906
rect 3903 10854 3917 10906
rect 3917 10854 3929 10906
rect 3929 10854 3959 10906
rect 3983 10854 3993 10906
rect 3993 10854 4039 10906
rect 3743 10852 3799 10854
rect 3823 10852 3879 10854
rect 3903 10852 3959 10854
rect 3983 10852 4039 10854
rect 3083 10362 3139 10364
rect 3163 10362 3219 10364
rect 3243 10362 3299 10364
rect 3323 10362 3379 10364
rect 3083 10310 3129 10362
rect 3129 10310 3139 10362
rect 3163 10310 3193 10362
rect 3193 10310 3205 10362
rect 3205 10310 3219 10362
rect 3243 10310 3257 10362
rect 3257 10310 3269 10362
rect 3269 10310 3299 10362
rect 3323 10310 3333 10362
rect 3333 10310 3379 10362
rect 3083 10308 3139 10310
rect 3163 10308 3219 10310
rect 3243 10308 3299 10310
rect 3323 10308 3379 10310
rect 3083 9274 3139 9276
rect 3163 9274 3219 9276
rect 3243 9274 3299 9276
rect 3323 9274 3379 9276
rect 3083 9222 3129 9274
rect 3129 9222 3139 9274
rect 3163 9222 3193 9274
rect 3193 9222 3205 9274
rect 3205 9222 3219 9274
rect 3243 9222 3257 9274
rect 3257 9222 3269 9274
rect 3269 9222 3299 9274
rect 3323 9222 3333 9274
rect 3333 9222 3379 9274
rect 3083 9220 3139 9222
rect 3163 9220 3219 9222
rect 3243 9220 3299 9222
rect 3323 9220 3379 9222
rect 3083 8186 3139 8188
rect 3163 8186 3219 8188
rect 3243 8186 3299 8188
rect 3323 8186 3379 8188
rect 3083 8134 3129 8186
rect 3129 8134 3139 8186
rect 3163 8134 3193 8186
rect 3193 8134 3205 8186
rect 3205 8134 3219 8186
rect 3243 8134 3257 8186
rect 3257 8134 3269 8186
rect 3269 8134 3299 8186
rect 3323 8134 3333 8186
rect 3333 8134 3379 8186
rect 3083 8132 3139 8134
rect 3163 8132 3219 8134
rect 3243 8132 3299 8134
rect 3323 8132 3379 8134
rect 3083 7098 3139 7100
rect 3163 7098 3219 7100
rect 3243 7098 3299 7100
rect 3323 7098 3379 7100
rect 3083 7046 3129 7098
rect 3129 7046 3139 7098
rect 3163 7046 3193 7098
rect 3193 7046 3205 7098
rect 3205 7046 3219 7098
rect 3243 7046 3257 7098
rect 3257 7046 3269 7098
rect 3269 7046 3299 7098
rect 3323 7046 3333 7098
rect 3333 7046 3379 7098
rect 3083 7044 3139 7046
rect 3163 7044 3219 7046
rect 3243 7044 3299 7046
rect 3323 7044 3379 7046
rect 3743 9818 3799 9820
rect 3823 9818 3879 9820
rect 3903 9818 3959 9820
rect 3983 9818 4039 9820
rect 3743 9766 3789 9818
rect 3789 9766 3799 9818
rect 3823 9766 3853 9818
rect 3853 9766 3865 9818
rect 3865 9766 3879 9818
rect 3903 9766 3917 9818
rect 3917 9766 3929 9818
rect 3929 9766 3959 9818
rect 3983 9766 3993 9818
rect 3993 9766 4039 9818
rect 3743 9764 3799 9766
rect 3823 9764 3879 9766
rect 3903 9764 3959 9766
rect 3983 9764 4039 9766
rect 4526 9560 4582 9616
rect 3743 8730 3799 8732
rect 3823 8730 3879 8732
rect 3903 8730 3959 8732
rect 3983 8730 4039 8732
rect 3743 8678 3789 8730
rect 3789 8678 3799 8730
rect 3823 8678 3853 8730
rect 3853 8678 3865 8730
rect 3865 8678 3879 8730
rect 3903 8678 3917 8730
rect 3917 8678 3929 8730
rect 3929 8678 3959 8730
rect 3983 8678 3993 8730
rect 3993 8678 4039 8730
rect 3743 8676 3799 8678
rect 3823 8676 3879 8678
rect 3903 8676 3959 8678
rect 3983 8676 4039 8678
rect 3606 8372 3608 8392
rect 3608 8372 3660 8392
rect 3660 8372 3662 8392
rect 3606 8336 3662 8372
rect 3743 7642 3799 7644
rect 3823 7642 3879 7644
rect 3903 7642 3959 7644
rect 3983 7642 4039 7644
rect 3743 7590 3789 7642
rect 3789 7590 3799 7642
rect 3823 7590 3853 7642
rect 3853 7590 3865 7642
rect 3865 7590 3879 7642
rect 3903 7590 3917 7642
rect 3917 7590 3929 7642
rect 3929 7590 3959 7642
rect 3983 7590 3993 7642
rect 3993 7590 4039 7642
rect 3743 7588 3799 7590
rect 3823 7588 3879 7590
rect 3903 7588 3959 7590
rect 3983 7588 4039 7590
rect 3743 6554 3799 6556
rect 3823 6554 3879 6556
rect 3903 6554 3959 6556
rect 3983 6554 4039 6556
rect 3743 6502 3789 6554
rect 3789 6502 3799 6554
rect 3823 6502 3853 6554
rect 3853 6502 3865 6554
rect 3865 6502 3879 6554
rect 3903 6502 3917 6554
rect 3917 6502 3929 6554
rect 3929 6502 3959 6554
rect 3983 6502 3993 6554
rect 3993 6502 4039 6554
rect 3743 6500 3799 6502
rect 3823 6500 3879 6502
rect 3903 6500 3959 6502
rect 3983 6500 4039 6502
rect 3083 6010 3139 6012
rect 3163 6010 3219 6012
rect 3243 6010 3299 6012
rect 3323 6010 3379 6012
rect 3083 5958 3129 6010
rect 3129 5958 3139 6010
rect 3163 5958 3193 6010
rect 3193 5958 3205 6010
rect 3205 5958 3219 6010
rect 3243 5958 3257 6010
rect 3257 5958 3269 6010
rect 3269 5958 3299 6010
rect 3323 5958 3333 6010
rect 3333 5958 3379 6010
rect 3083 5956 3139 5958
rect 3163 5956 3219 5958
rect 3243 5956 3299 5958
rect 3323 5956 3379 5958
rect 3083 4922 3139 4924
rect 3163 4922 3219 4924
rect 3243 4922 3299 4924
rect 3323 4922 3379 4924
rect 3083 4870 3129 4922
rect 3129 4870 3139 4922
rect 3163 4870 3193 4922
rect 3193 4870 3205 4922
rect 3205 4870 3219 4922
rect 3243 4870 3257 4922
rect 3257 4870 3269 4922
rect 3269 4870 3299 4922
rect 3323 4870 3333 4922
rect 3333 4870 3379 4922
rect 3083 4868 3139 4870
rect 3163 4868 3219 4870
rect 3243 4868 3299 4870
rect 3323 4868 3379 4870
rect 3743 5466 3799 5468
rect 3823 5466 3879 5468
rect 3903 5466 3959 5468
rect 3983 5466 4039 5468
rect 3743 5414 3789 5466
rect 3789 5414 3799 5466
rect 3823 5414 3853 5466
rect 3853 5414 3865 5466
rect 3865 5414 3879 5466
rect 3903 5414 3917 5466
rect 3917 5414 3929 5466
rect 3929 5414 3959 5466
rect 3983 5414 3993 5466
rect 3993 5414 4039 5466
rect 3743 5412 3799 5414
rect 3823 5412 3879 5414
rect 3903 5412 3959 5414
rect 3983 5412 4039 5414
rect 4434 6840 4490 6896
rect 5998 13368 6054 13424
rect 11593 19066 11649 19068
rect 11673 19066 11729 19068
rect 11753 19066 11809 19068
rect 11833 19066 11889 19068
rect 11593 19014 11639 19066
rect 11639 19014 11649 19066
rect 11673 19014 11703 19066
rect 11703 19014 11715 19066
rect 11715 19014 11729 19066
rect 11753 19014 11767 19066
rect 11767 19014 11779 19066
rect 11779 19014 11809 19066
rect 11833 19014 11843 19066
rect 11843 19014 11889 19066
rect 11593 19012 11649 19014
rect 11673 19012 11729 19014
rect 11753 19012 11809 19014
rect 11833 19012 11889 19014
rect 15848 19066 15904 19068
rect 15928 19066 15984 19068
rect 16008 19066 16064 19068
rect 16088 19066 16144 19068
rect 15848 19014 15894 19066
rect 15894 19014 15904 19066
rect 15928 19014 15958 19066
rect 15958 19014 15970 19066
rect 15970 19014 15984 19066
rect 16008 19014 16022 19066
rect 16022 19014 16034 19066
rect 16034 19014 16064 19066
rect 16088 19014 16098 19066
rect 16098 19014 16144 19066
rect 15848 19012 15904 19014
rect 15928 19012 15984 19014
rect 16008 19012 16064 19014
rect 16088 19012 16144 19014
rect 7998 16346 8054 16348
rect 8078 16346 8134 16348
rect 8158 16346 8214 16348
rect 8238 16346 8294 16348
rect 7998 16294 8044 16346
rect 8044 16294 8054 16346
rect 8078 16294 8108 16346
rect 8108 16294 8120 16346
rect 8120 16294 8134 16346
rect 8158 16294 8172 16346
rect 8172 16294 8184 16346
rect 8184 16294 8214 16346
rect 8238 16294 8248 16346
rect 8248 16294 8294 16346
rect 7998 16292 8054 16294
rect 8078 16292 8134 16294
rect 8158 16292 8214 16294
rect 8238 16292 8294 16294
rect 7338 15802 7394 15804
rect 7418 15802 7474 15804
rect 7498 15802 7554 15804
rect 7578 15802 7634 15804
rect 7338 15750 7384 15802
rect 7384 15750 7394 15802
rect 7418 15750 7448 15802
rect 7448 15750 7460 15802
rect 7460 15750 7474 15802
rect 7498 15750 7512 15802
rect 7512 15750 7524 15802
rect 7524 15750 7554 15802
rect 7578 15750 7588 15802
rect 7588 15750 7634 15802
rect 7338 15748 7394 15750
rect 7418 15748 7474 15750
rect 7498 15748 7554 15750
rect 7578 15748 7634 15750
rect 4894 6704 4950 6760
rect 3743 4378 3799 4380
rect 3823 4378 3879 4380
rect 3903 4378 3959 4380
rect 3983 4378 4039 4380
rect 3743 4326 3789 4378
rect 3789 4326 3799 4378
rect 3823 4326 3853 4378
rect 3853 4326 3865 4378
rect 3865 4326 3879 4378
rect 3903 4326 3917 4378
rect 3917 4326 3929 4378
rect 3929 4326 3959 4378
rect 3983 4326 3993 4378
rect 3993 4326 4039 4378
rect 3743 4324 3799 4326
rect 3823 4324 3879 4326
rect 3903 4324 3959 4326
rect 3983 4324 4039 4326
rect 3083 3834 3139 3836
rect 3163 3834 3219 3836
rect 3243 3834 3299 3836
rect 3323 3834 3379 3836
rect 3083 3782 3129 3834
rect 3129 3782 3139 3834
rect 3163 3782 3193 3834
rect 3193 3782 3205 3834
rect 3205 3782 3219 3834
rect 3243 3782 3257 3834
rect 3257 3782 3269 3834
rect 3269 3782 3299 3834
rect 3323 3782 3333 3834
rect 3333 3782 3379 3834
rect 3083 3780 3139 3782
rect 3163 3780 3219 3782
rect 3243 3780 3299 3782
rect 3323 3780 3379 3782
rect 5354 5072 5410 5128
rect 5170 4684 5226 4720
rect 5170 4664 5172 4684
rect 5172 4664 5224 4684
rect 5224 4664 5226 4684
rect 6090 6568 6146 6624
rect 6182 6196 6184 6216
rect 6184 6196 6236 6216
rect 6236 6196 6238 6216
rect 6182 6160 6238 6196
rect 7338 14714 7394 14716
rect 7418 14714 7474 14716
rect 7498 14714 7554 14716
rect 7578 14714 7634 14716
rect 7338 14662 7384 14714
rect 7384 14662 7394 14714
rect 7418 14662 7448 14714
rect 7448 14662 7460 14714
rect 7460 14662 7474 14714
rect 7498 14662 7512 14714
rect 7512 14662 7524 14714
rect 7524 14662 7554 14714
rect 7578 14662 7588 14714
rect 7588 14662 7634 14714
rect 7338 14660 7394 14662
rect 7418 14660 7474 14662
rect 7498 14660 7554 14662
rect 7578 14660 7634 14662
rect 7998 15258 8054 15260
rect 8078 15258 8134 15260
rect 8158 15258 8214 15260
rect 8238 15258 8294 15260
rect 7998 15206 8044 15258
rect 8044 15206 8054 15258
rect 8078 15206 8108 15258
rect 8108 15206 8120 15258
rect 8120 15206 8134 15258
rect 8158 15206 8172 15258
rect 8172 15206 8184 15258
rect 8184 15206 8214 15258
rect 8238 15206 8248 15258
rect 8248 15206 8294 15258
rect 7998 15204 8054 15206
rect 8078 15204 8134 15206
rect 8158 15204 8214 15206
rect 8238 15204 8294 15206
rect 7998 14170 8054 14172
rect 8078 14170 8134 14172
rect 8158 14170 8214 14172
rect 8238 14170 8294 14172
rect 7998 14118 8044 14170
rect 8044 14118 8054 14170
rect 8078 14118 8108 14170
rect 8108 14118 8120 14170
rect 8120 14118 8134 14170
rect 8158 14118 8172 14170
rect 8172 14118 8184 14170
rect 8184 14118 8214 14170
rect 8238 14118 8248 14170
rect 8248 14118 8294 14170
rect 7998 14116 8054 14118
rect 8078 14116 8134 14118
rect 8158 14116 8214 14118
rect 8238 14116 8294 14118
rect 7338 13626 7394 13628
rect 7418 13626 7474 13628
rect 7498 13626 7554 13628
rect 7578 13626 7634 13628
rect 7338 13574 7384 13626
rect 7384 13574 7394 13626
rect 7418 13574 7448 13626
rect 7448 13574 7460 13626
rect 7460 13574 7474 13626
rect 7498 13574 7512 13626
rect 7512 13574 7524 13626
rect 7524 13574 7554 13626
rect 7578 13574 7588 13626
rect 7588 13574 7634 13626
rect 7338 13572 7394 13574
rect 7418 13572 7474 13574
rect 7498 13572 7554 13574
rect 7578 13572 7634 13574
rect 7338 12538 7394 12540
rect 7418 12538 7474 12540
rect 7498 12538 7554 12540
rect 7578 12538 7634 12540
rect 7338 12486 7384 12538
rect 7384 12486 7394 12538
rect 7418 12486 7448 12538
rect 7448 12486 7460 12538
rect 7460 12486 7474 12538
rect 7498 12486 7512 12538
rect 7512 12486 7524 12538
rect 7524 12486 7554 12538
rect 7578 12486 7588 12538
rect 7588 12486 7634 12538
rect 7338 12484 7394 12486
rect 7418 12484 7474 12486
rect 7498 12484 7554 12486
rect 7578 12484 7634 12486
rect 7338 11450 7394 11452
rect 7418 11450 7474 11452
rect 7498 11450 7554 11452
rect 7578 11450 7634 11452
rect 7338 11398 7384 11450
rect 7384 11398 7394 11450
rect 7418 11398 7448 11450
rect 7448 11398 7460 11450
rect 7460 11398 7474 11450
rect 7498 11398 7512 11450
rect 7512 11398 7524 11450
rect 7524 11398 7554 11450
rect 7578 11398 7588 11450
rect 7588 11398 7634 11450
rect 7338 11396 7394 11398
rect 7418 11396 7474 11398
rect 7498 11396 7554 11398
rect 7578 11396 7634 11398
rect 3743 3290 3799 3292
rect 3823 3290 3879 3292
rect 3903 3290 3959 3292
rect 3983 3290 4039 3292
rect 3743 3238 3789 3290
rect 3789 3238 3799 3290
rect 3823 3238 3853 3290
rect 3853 3238 3865 3290
rect 3865 3238 3879 3290
rect 3903 3238 3917 3290
rect 3917 3238 3929 3290
rect 3929 3238 3959 3290
rect 3983 3238 3993 3290
rect 3993 3238 4039 3290
rect 3743 3236 3799 3238
rect 3823 3236 3879 3238
rect 3903 3236 3959 3238
rect 3983 3236 4039 3238
rect 3083 2746 3139 2748
rect 3163 2746 3219 2748
rect 3243 2746 3299 2748
rect 3323 2746 3379 2748
rect 3083 2694 3129 2746
rect 3129 2694 3139 2746
rect 3163 2694 3193 2746
rect 3193 2694 3205 2746
rect 3205 2694 3219 2746
rect 3243 2694 3257 2746
rect 3257 2694 3269 2746
rect 3269 2694 3299 2746
rect 3323 2694 3333 2746
rect 3333 2694 3379 2746
rect 3083 2692 3139 2694
rect 3163 2692 3219 2694
rect 3243 2692 3299 2694
rect 3323 2692 3379 2694
rect 7338 10362 7394 10364
rect 7418 10362 7474 10364
rect 7498 10362 7554 10364
rect 7578 10362 7634 10364
rect 7338 10310 7384 10362
rect 7384 10310 7394 10362
rect 7418 10310 7448 10362
rect 7448 10310 7460 10362
rect 7460 10310 7474 10362
rect 7498 10310 7512 10362
rect 7512 10310 7524 10362
rect 7524 10310 7554 10362
rect 7578 10310 7588 10362
rect 7588 10310 7634 10362
rect 7338 10308 7394 10310
rect 7418 10308 7474 10310
rect 7498 10308 7554 10310
rect 7578 10308 7634 10310
rect 7998 13082 8054 13084
rect 8078 13082 8134 13084
rect 8158 13082 8214 13084
rect 8238 13082 8294 13084
rect 7998 13030 8044 13082
rect 8044 13030 8054 13082
rect 8078 13030 8108 13082
rect 8108 13030 8120 13082
rect 8120 13030 8134 13082
rect 8158 13030 8172 13082
rect 8172 13030 8184 13082
rect 8184 13030 8214 13082
rect 8238 13030 8248 13082
rect 8248 13030 8294 13082
rect 7998 13028 8054 13030
rect 8078 13028 8134 13030
rect 8158 13028 8214 13030
rect 8238 13028 8294 13030
rect 12253 18522 12309 18524
rect 12333 18522 12389 18524
rect 12413 18522 12469 18524
rect 12493 18522 12549 18524
rect 12253 18470 12299 18522
rect 12299 18470 12309 18522
rect 12333 18470 12363 18522
rect 12363 18470 12375 18522
rect 12375 18470 12389 18522
rect 12413 18470 12427 18522
rect 12427 18470 12439 18522
rect 12439 18470 12469 18522
rect 12493 18470 12503 18522
rect 12503 18470 12549 18522
rect 12253 18468 12309 18470
rect 12333 18468 12389 18470
rect 12413 18468 12469 18470
rect 12493 18468 12549 18470
rect 11593 17978 11649 17980
rect 11673 17978 11729 17980
rect 11753 17978 11809 17980
rect 11833 17978 11889 17980
rect 11593 17926 11639 17978
rect 11639 17926 11649 17978
rect 11673 17926 11703 17978
rect 11703 17926 11715 17978
rect 11715 17926 11729 17978
rect 11753 17926 11767 17978
rect 11767 17926 11779 17978
rect 11779 17926 11809 17978
rect 11833 17926 11843 17978
rect 11843 17926 11889 17978
rect 11593 17924 11649 17926
rect 11673 17924 11729 17926
rect 11753 17924 11809 17926
rect 11833 17924 11889 17926
rect 8758 13776 8814 13832
rect 7998 11994 8054 11996
rect 8078 11994 8134 11996
rect 8158 11994 8214 11996
rect 8238 11994 8294 11996
rect 7998 11942 8044 11994
rect 8044 11942 8054 11994
rect 8078 11942 8108 11994
rect 8108 11942 8120 11994
rect 8120 11942 8134 11994
rect 8158 11942 8172 11994
rect 8172 11942 8184 11994
rect 8184 11942 8214 11994
rect 8238 11942 8248 11994
rect 8248 11942 8294 11994
rect 7998 11940 8054 11942
rect 8078 11940 8134 11942
rect 8158 11940 8214 11942
rect 8238 11940 8294 11942
rect 7998 10906 8054 10908
rect 8078 10906 8134 10908
rect 8158 10906 8214 10908
rect 8238 10906 8294 10908
rect 7998 10854 8044 10906
rect 8044 10854 8054 10906
rect 8078 10854 8108 10906
rect 8108 10854 8120 10906
rect 8120 10854 8134 10906
rect 8158 10854 8172 10906
rect 8172 10854 8184 10906
rect 8184 10854 8214 10906
rect 8238 10854 8248 10906
rect 8248 10854 8294 10906
rect 7998 10852 8054 10854
rect 8078 10852 8134 10854
rect 8158 10852 8214 10854
rect 8238 10852 8294 10854
rect 7338 9274 7394 9276
rect 7418 9274 7474 9276
rect 7498 9274 7554 9276
rect 7578 9274 7634 9276
rect 7338 9222 7384 9274
rect 7384 9222 7394 9274
rect 7418 9222 7448 9274
rect 7448 9222 7460 9274
rect 7460 9222 7474 9274
rect 7498 9222 7512 9274
rect 7512 9222 7524 9274
rect 7524 9222 7554 9274
rect 7578 9222 7588 9274
rect 7588 9222 7634 9274
rect 7338 9220 7394 9222
rect 7418 9220 7474 9222
rect 7498 9220 7554 9222
rect 7578 9220 7634 9222
rect 7998 9818 8054 9820
rect 8078 9818 8134 9820
rect 8158 9818 8214 9820
rect 8238 9818 8294 9820
rect 7998 9766 8044 9818
rect 8044 9766 8054 9818
rect 8078 9766 8108 9818
rect 8108 9766 8120 9818
rect 8120 9766 8134 9818
rect 8158 9766 8172 9818
rect 8172 9766 8184 9818
rect 8184 9766 8214 9818
rect 8238 9766 8248 9818
rect 8248 9766 8294 9818
rect 7998 9764 8054 9766
rect 8078 9764 8134 9766
rect 8158 9764 8214 9766
rect 8238 9764 8294 9766
rect 6918 5616 6974 5672
rect 6550 4820 6606 4856
rect 6550 4800 6552 4820
rect 6552 4800 6604 4820
rect 6604 4800 6606 4820
rect 7010 5092 7066 5128
rect 7010 5072 7012 5092
rect 7012 5072 7064 5092
rect 7064 5072 7066 5092
rect 6918 4800 6974 4856
rect 6826 4528 6882 4584
rect 7338 8186 7394 8188
rect 7418 8186 7474 8188
rect 7498 8186 7554 8188
rect 7578 8186 7634 8188
rect 7338 8134 7384 8186
rect 7384 8134 7394 8186
rect 7418 8134 7448 8186
rect 7448 8134 7460 8186
rect 7460 8134 7474 8186
rect 7498 8134 7512 8186
rect 7512 8134 7524 8186
rect 7524 8134 7554 8186
rect 7578 8134 7588 8186
rect 7588 8134 7634 8186
rect 7338 8132 7394 8134
rect 7418 8132 7474 8134
rect 7498 8132 7554 8134
rect 7578 8132 7634 8134
rect 7378 7928 7434 7984
rect 7338 7098 7394 7100
rect 7418 7098 7474 7100
rect 7498 7098 7554 7100
rect 7578 7098 7634 7100
rect 7338 7046 7384 7098
rect 7384 7046 7394 7098
rect 7418 7046 7448 7098
rect 7448 7046 7460 7098
rect 7460 7046 7474 7098
rect 7498 7046 7512 7098
rect 7512 7046 7524 7098
rect 7524 7046 7554 7098
rect 7578 7046 7588 7098
rect 7588 7046 7634 7098
rect 7338 7044 7394 7046
rect 7418 7044 7474 7046
rect 7498 7044 7554 7046
rect 7578 7044 7634 7046
rect 7378 6568 7434 6624
rect 7286 6160 7342 6216
rect 7338 6010 7394 6012
rect 7418 6010 7474 6012
rect 7498 6010 7554 6012
rect 7578 6010 7634 6012
rect 7338 5958 7384 6010
rect 7384 5958 7394 6010
rect 7418 5958 7448 6010
rect 7448 5958 7460 6010
rect 7460 5958 7474 6010
rect 7498 5958 7512 6010
rect 7512 5958 7524 6010
rect 7524 5958 7554 6010
rect 7578 5958 7588 6010
rect 7588 5958 7634 6010
rect 7338 5956 7394 5958
rect 7418 5956 7474 5958
rect 7498 5956 7554 5958
rect 7578 5956 7634 5958
rect 7194 5616 7250 5672
rect 7998 8730 8054 8732
rect 8078 8730 8134 8732
rect 8158 8730 8214 8732
rect 8238 8730 8294 8732
rect 7998 8678 8044 8730
rect 8044 8678 8054 8730
rect 8078 8678 8108 8730
rect 8108 8678 8120 8730
rect 8120 8678 8134 8730
rect 8158 8678 8172 8730
rect 8172 8678 8184 8730
rect 8184 8678 8214 8730
rect 8238 8678 8248 8730
rect 8248 8678 8294 8730
rect 7998 8676 8054 8678
rect 8078 8676 8134 8678
rect 8158 8676 8214 8678
rect 8238 8676 8294 8678
rect 7998 7642 8054 7644
rect 8078 7642 8134 7644
rect 8158 7642 8214 7644
rect 8238 7642 8294 7644
rect 7998 7590 8044 7642
rect 8044 7590 8054 7642
rect 8078 7590 8108 7642
rect 8108 7590 8120 7642
rect 8120 7590 8134 7642
rect 8158 7590 8172 7642
rect 8172 7590 8184 7642
rect 8184 7590 8214 7642
rect 8238 7590 8248 7642
rect 8248 7590 8294 7642
rect 7998 7588 8054 7590
rect 8078 7588 8134 7590
rect 8158 7588 8214 7590
rect 8238 7588 8294 7590
rect 7998 6554 8054 6556
rect 8078 6554 8134 6556
rect 8158 6554 8214 6556
rect 8238 6554 8294 6556
rect 7998 6502 8044 6554
rect 8044 6502 8054 6554
rect 8078 6502 8108 6554
rect 8108 6502 8120 6554
rect 8120 6502 8134 6554
rect 8158 6502 8172 6554
rect 8172 6502 8184 6554
rect 8184 6502 8214 6554
rect 8238 6502 8248 6554
rect 8248 6502 8294 6554
rect 7998 6500 8054 6502
rect 8078 6500 8134 6502
rect 8158 6500 8214 6502
rect 8238 6500 8294 6502
rect 7338 4922 7394 4924
rect 7418 4922 7474 4924
rect 7498 4922 7554 4924
rect 7578 4922 7634 4924
rect 7338 4870 7384 4922
rect 7384 4870 7394 4922
rect 7418 4870 7448 4922
rect 7448 4870 7460 4922
rect 7460 4870 7474 4922
rect 7498 4870 7512 4922
rect 7512 4870 7524 4922
rect 7524 4870 7554 4922
rect 7578 4870 7588 4922
rect 7588 4870 7634 4922
rect 7338 4868 7394 4870
rect 7418 4868 7474 4870
rect 7498 4868 7554 4870
rect 7578 4868 7634 4870
rect 7286 4564 7288 4584
rect 7288 4564 7340 4584
rect 7340 4564 7342 4584
rect 7286 4528 7342 4564
rect 7338 3834 7394 3836
rect 7418 3834 7474 3836
rect 7498 3834 7554 3836
rect 7578 3834 7634 3836
rect 7338 3782 7384 3834
rect 7384 3782 7394 3834
rect 7418 3782 7448 3834
rect 7448 3782 7460 3834
rect 7460 3782 7474 3834
rect 7498 3782 7512 3834
rect 7512 3782 7524 3834
rect 7524 3782 7554 3834
rect 7578 3782 7588 3834
rect 7588 3782 7634 3834
rect 7338 3780 7394 3782
rect 7418 3780 7474 3782
rect 7498 3780 7554 3782
rect 7578 3780 7634 3782
rect 7338 2746 7394 2748
rect 7418 2746 7474 2748
rect 7498 2746 7554 2748
rect 7578 2746 7634 2748
rect 7338 2694 7384 2746
rect 7384 2694 7394 2746
rect 7418 2694 7448 2746
rect 7448 2694 7460 2746
rect 7460 2694 7474 2746
rect 7498 2694 7512 2746
rect 7512 2694 7524 2746
rect 7524 2694 7554 2746
rect 7578 2694 7588 2746
rect 7588 2694 7634 2746
rect 7338 2692 7394 2694
rect 7418 2692 7474 2694
rect 7498 2692 7554 2694
rect 7578 2692 7634 2694
rect 7998 5466 8054 5468
rect 8078 5466 8134 5468
rect 8158 5466 8214 5468
rect 8238 5466 8294 5468
rect 7998 5414 8044 5466
rect 8044 5414 8054 5466
rect 8078 5414 8108 5466
rect 8108 5414 8120 5466
rect 8120 5414 8134 5466
rect 8158 5414 8172 5466
rect 8172 5414 8184 5466
rect 8184 5414 8214 5466
rect 8238 5414 8248 5466
rect 8248 5414 8294 5466
rect 7998 5412 8054 5414
rect 8078 5412 8134 5414
rect 8158 5412 8214 5414
rect 8238 5412 8294 5414
rect 8022 5092 8078 5128
rect 8022 5072 8024 5092
rect 8024 5072 8076 5092
rect 8076 5072 8078 5092
rect 7998 4378 8054 4380
rect 8078 4378 8134 4380
rect 8158 4378 8214 4380
rect 8238 4378 8294 4380
rect 7998 4326 8044 4378
rect 8044 4326 8054 4378
rect 8078 4326 8108 4378
rect 8108 4326 8120 4378
rect 8120 4326 8134 4378
rect 8158 4326 8172 4378
rect 8172 4326 8184 4378
rect 8184 4326 8214 4378
rect 8238 4326 8248 4378
rect 8248 4326 8294 4378
rect 7998 4324 8054 4326
rect 8078 4324 8134 4326
rect 8158 4324 8214 4326
rect 8238 4324 8294 4326
rect 7998 3290 8054 3292
rect 8078 3290 8134 3292
rect 8158 3290 8214 3292
rect 8238 3290 8294 3292
rect 7998 3238 8044 3290
rect 8044 3238 8054 3290
rect 8078 3238 8108 3290
rect 8108 3238 8120 3290
rect 8120 3238 8134 3290
rect 8158 3238 8172 3290
rect 8172 3238 8184 3290
rect 8184 3238 8214 3290
rect 8238 3238 8248 3290
rect 8248 3238 8294 3290
rect 7998 3236 8054 3238
rect 8078 3236 8134 3238
rect 8158 3236 8214 3238
rect 8238 3236 8294 3238
rect 9494 10668 9550 10704
rect 9494 10648 9496 10668
rect 9496 10648 9548 10668
rect 9548 10648 9550 10668
rect 9034 4664 9090 4720
rect 3743 2202 3799 2204
rect 3823 2202 3879 2204
rect 3903 2202 3959 2204
rect 3983 2202 4039 2204
rect 3743 2150 3789 2202
rect 3789 2150 3799 2202
rect 3823 2150 3853 2202
rect 3853 2150 3865 2202
rect 3865 2150 3879 2202
rect 3903 2150 3917 2202
rect 3917 2150 3929 2202
rect 3929 2150 3959 2202
rect 3983 2150 3993 2202
rect 3993 2150 4039 2202
rect 3743 2148 3799 2150
rect 3823 2148 3879 2150
rect 3903 2148 3959 2150
rect 3983 2148 4039 2150
rect 7998 2202 8054 2204
rect 8078 2202 8134 2204
rect 8158 2202 8214 2204
rect 8238 2202 8294 2204
rect 7998 2150 8044 2202
rect 8044 2150 8054 2202
rect 8078 2150 8108 2202
rect 8108 2150 8120 2202
rect 8120 2150 8134 2202
rect 8158 2150 8172 2202
rect 8172 2150 8184 2202
rect 8184 2150 8214 2202
rect 8238 2150 8248 2202
rect 8248 2150 8294 2202
rect 7998 2148 8054 2150
rect 8078 2148 8134 2150
rect 8158 2148 8214 2150
rect 8238 2148 8294 2150
rect 9494 6840 9550 6896
rect 9954 6840 10010 6896
rect 10782 10804 10838 10840
rect 10782 10784 10784 10804
rect 10784 10784 10836 10804
rect 10836 10784 10838 10804
rect 10690 9560 10746 9616
rect 11593 16890 11649 16892
rect 11673 16890 11729 16892
rect 11753 16890 11809 16892
rect 11833 16890 11889 16892
rect 11593 16838 11639 16890
rect 11639 16838 11649 16890
rect 11673 16838 11703 16890
rect 11703 16838 11715 16890
rect 11715 16838 11729 16890
rect 11753 16838 11767 16890
rect 11767 16838 11779 16890
rect 11779 16838 11809 16890
rect 11833 16838 11843 16890
rect 11843 16838 11889 16890
rect 11593 16836 11649 16838
rect 11673 16836 11729 16838
rect 11753 16836 11809 16838
rect 11833 16836 11889 16838
rect 12253 17434 12309 17436
rect 12333 17434 12389 17436
rect 12413 17434 12469 17436
rect 12493 17434 12549 17436
rect 12253 17382 12299 17434
rect 12299 17382 12309 17434
rect 12333 17382 12363 17434
rect 12363 17382 12375 17434
rect 12375 17382 12389 17434
rect 12413 17382 12427 17434
rect 12427 17382 12439 17434
rect 12439 17382 12469 17434
rect 12493 17382 12503 17434
rect 12503 17382 12549 17434
rect 12253 17380 12309 17382
rect 12333 17380 12389 17382
rect 12413 17380 12469 17382
rect 12493 17380 12549 17382
rect 12253 16346 12309 16348
rect 12333 16346 12389 16348
rect 12413 16346 12469 16348
rect 12493 16346 12549 16348
rect 12253 16294 12299 16346
rect 12299 16294 12309 16346
rect 12333 16294 12363 16346
rect 12363 16294 12375 16346
rect 12375 16294 12389 16346
rect 12413 16294 12427 16346
rect 12427 16294 12439 16346
rect 12439 16294 12469 16346
rect 12493 16294 12503 16346
rect 12503 16294 12549 16346
rect 12253 16292 12309 16294
rect 12333 16292 12389 16294
rect 12413 16292 12469 16294
rect 12493 16292 12549 16294
rect 11593 15802 11649 15804
rect 11673 15802 11729 15804
rect 11753 15802 11809 15804
rect 11833 15802 11889 15804
rect 11593 15750 11639 15802
rect 11639 15750 11649 15802
rect 11673 15750 11703 15802
rect 11703 15750 11715 15802
rect 11715 15750 11729 15802
rect 11753 15750 11767 15802
rect 11767 15750 11779 15802
rect 11779 15750 11809 15802
rect 11833 15750 11843 15802
rect 11843 15750 11889 15802
rect 11593 15748 11649 15750
rect 11673 15748 11729 15750
rect 11753 15748 11809 15750
rect 11833 15748 11889 15750
rect 12253 15258 12309 15260
rect 12333 15258 12389 15260
rect 12413 15258 12469 15260
rect 12493 15258 12549 15260
rect 12253 15206 12299 15258
rect 12299 15206 12309 15258
rect 12333 15206 12363 15258
rect 12363 15206 12375 15258
rect 12375 15206 12389 15258
rect 12413 15206 12427 15258
rect 12427 15206 12439 15258
rect 12439 15206 12469 15258
rect 12493 15206 12503 15258
rect 12503 15206 12549 15258
rect 12253 15204 12309 15206
rect 12333 15204 12389 15206
rect 12413 15204 12469 15206
rect 12493 15204 12549 15206
rect 11593 14714 11649 14716
rect 11673 14714 11729 14716
rect 11753 14714 11809 14716
rect 11833 14714 11889 14716
rect 11593 14662 11639 14714
rect 11639 14662 11649 14714
rect 11673 14662 11703 14714
rect 11703 14662 11715 14714
rect 11715 14662 11729 14714
rect 11753 14662 11767 14714
rect 11767 14662 11779 14714
rect 11779 14662 11809 14714
rect 11833 14662 11843 14714
rect 11843 14662 11889 14714
rect 11593 14660 11649 14662
rect 11673 14660 11729 14662
rect 11753 14660 11809 14662
rect 11833 14660 11889 14662
rect 12253 14170 12309 14172
rect 12333 14170 12389 14172
rect 12413 14170 12469 14172
rect 12493 14170 12549 14172
rect 12253 14118 12299 14170
rect 12299 14118 12309 14170
rect 12333 14118 12363 14170
rect 12363 14118 12375 14170
rect 12375 14118 12389 14170
rect 12413 14118 12427 14170
rect 12427 14118 12439 14170
rect 12439 14118 12469 14170
rect 12493 14118 12503 14170
rect 12503 14118 12549 14170
rect 12253 14116 12309 14118
rect 12333 14116 12389 14118
rect 12413 14116 12469 14118
rect 12493 14116 12549 14118
rect 12714 15000 12770 15056
rect 11593 13626 11649 13628
rect 11673 13626 11729 13628
rect 11753 13626 11809 13628
rect 11833 13626 11889 13628
rect 11593 13574 11639 13626
rect 11639 13574 11649 13626
rect 11673 13574 11703 13626
rect 11703 13574 11715 13626
rect 11715 13574 11729 13626
rect 11753 13574 11767 13626
rect 11767 13574 11779 13626
rect 11779 13574 11809 13626
rect 11833 13574 11843 13626
rect 11843 13574 11889 13626
rect 11593 13572 11649 13574
rect 11673 13572 11729 13574
rect 11753 13572 11809 13574
rect 11833 13572 11889 13574
rect 12253 13082 12309 13084
rect 12333 13082 12389 13084
rect 12413 13082 12469 13084
rect 12493 13082 12549 13084
rect 12253 13030 12299 13082
rect 12299 13030 12309 13082
rect 12333 13030 12363 13082
rect 12363 13030 12375 13082
rect 12375 13030 12389 13082
rect 12413 13030 12427 13082
rect 12427 13030 12439 13082
rect 12439 13030 12469 13082
rect 12493 13030 12503 13082
rect 12503 13030 12549 13082
rect 12253 13028 12309 13030
rect 12333 13028 12389 13030
rect 12413 13028 12469 13030
rect 12493 13028 12549 13030
rect 11593 12538 11649 12540
rect 11673 12538 11729 12540
rect 11753 12538 11809 12540
rect 11833 12538 11889 12540
rect 11593 12486 11639 12538
rect 11639 12486 11649 12538
rect 11673 12486 11703 12538
rect 11703 12486 11715 12538
rect 11715 12486 11729 12538
rect 11753 12486 11767 12538
rect 11767 12486 11779 12538
rect 11779 12486 11809 12538
rect 11833 12486 11843 12538
rect 11843 12486 11889 12538
rect 11593 12484 11649 12486
rect 11673 12484 11729 12486
rect 11753 12484 11809 12486
rect 11833 12484 11889 12486
rect 12253 11994 12309 11996
rect 12333 11994 12389 11996
rect 12413 11994 12469 11996
rect 12493 11994 12549 11996
rect 12253 11942 12299 11994
rect 12299 11942 12309 11994
rect 12333 11942 12363 11994
rect 12363 11942 12375 11994
rect 12375 11942 12389 11994
rect 12413 11942 12427 11994
rect 12427 11942 12439 11994
rect 12439 11942 12469 11994
rect 12493 11942 12503 11994
rect 12503 11942 12549 11994
rect 12253 11940 12309 11942
rect 12333 11940 12389 11942
rect 12413 11940 12469 11942
rect 12493 11940 12549 11942
rect 11593 11450 11649 11452
rect 11673 11450 11729 11452
rect 11753 11450 11809 11452
rect 11833 11450 11889 11452
rect 11593 11398 11639 11450
rect 11639 11398 11649 11450
rect 11673 11398 11703 11450
rect 11703 11398 11715 11450
rect 11715 11398 11729 11450
rect 11753 11398 11767 11450
rect 11767 11398 11779 11450
rect 11779 11398 11809 11450
rect 11833 11398 11843 11450
rect 11843 11398 11889 11450
rect 11593 11396 11649 11398
rect 11673 11396 11729 11398
rect 11753 11396 11809 11398
rect 11833 11396 11889 11398
rect 12253 10906 12309 10908
rect 12333 10906 12389 10908
rect 12413 10906 12469 10908
rect 12493 10906 12549 10908
rect 12253 10854 12299 10906
rect 12299 10854 12309 10906
rect 12333 10854 12363 10906
rect 12363 10854 12375 10906
rect 12375 10854 12389 10906
rect 12413 10854 12427 10906
rect 12427 10854 12439 10906
rect 12439 10854 12469 10906
rect 12493 10854 12503 10906
rect 12503 10854 12549 10906
rect 12253 10852 12309 10854
rect 12333 10852 12389 10854
rect 12413 10852 12469 10854
rect 12493 10852 12549 10854
rect 11593 10362 11649 10364
rect 11673 10362 11729 10364
rect 11753 10362 11809 10364
rect 11833 10362 11889 10364
rect 11593 10310 11639 10362
rect 11639 10310 11649 10362
rect 11673 10310 11703 10362
rect 11703 10310 11715 10362
rect 11715 10310 11729 10362
rect 11753 10310 11767 10362
rect 11767 10310 11779 10362
rect 11779 10310 11809 10362
rect 11833 10310 11843 10362
rect 11843 10310 11889 10362
rect 11593 10308 11649 10310
rect 11673 10308 11729 10310
rect 11753 10308 11809 10310
rect 11833 10308 11889 10310
rect 11702 9560 11758 9616
rect 11593 9274 11649 9276
rect 11673 9274 11729 9276
rect 11753 9274 11809 9276
rect 11833 9274 11889 9276
rect 11593 9222 11639 9274
rect 11639 9222 11649 9274
rect 11673 9222 11703 9274
rect 11703 9222 11715 9274
rect 11715 9222 11729 9274
rect 11753 9222 11767 9274
rect 11767 9222 11779 9274
rect 11779 9222 11809 9274
rect 11833 9222 11843 9274
rect 11843 9222 11889 9274
rect 11593 9220 11649 9222
rect 11673 9220 11729 9222
rect 11753 9220 11809 9222
rect 11833 9220 11889 9222
rect 11242 8336 11298 8392
rect 10138 2896 10194 2952
rect 11593 8186 11649 8188
rect 11673 8186 11729 8188
rect 11753 8186 11809 8188
rect 11833 8186 11889 8188
rect 11593 8134 11639 8186
rect 11639 8134 11649 8186
rect 11673 8134 11703 8186
rect 11703 8134 11715 8186
rect 11715 8134 11729 8186
rect 11753 8134 11767 8186
rect 11767 8134 11779 8186
rect 11779 8134 11809 8186
rect 11833 8134 11843 8186
rect 11843 8134 11889 8186
rect 11593 8132 11649 8134
rect 11673 8132 11729 8134
rect 11753 8132 11809 8134
rect 11833 8132 11889 8134
rect 12253 9818 12309 9820
rect 12333 9818 12389 9820
rect 12413 9818 12469 9820
rect 12493 9818 12549 9820
rect 12253 9766 12299 9818
rect 12299 9766 12309 9818
rect 12333 9766 12363 9818
rect 12363 9766 12375 9818
rect 12375 9766 12389 9818
rect 12413 9766 12427 9818
rect 12427 9766 12439 9818
rect 12439 9766 12469 9818
rect 12493 9766 12503 9818
rect 12503 9766 12549 9818
rect 12253 9764 12309 9766
rect 12333 9764 12389 9766
rect 12413 9764 12469 9766
rect 12493 9764 12549 9766
rect 12253 8730 12309 8732
rect 12333 8730 12389 8732
rect 12413 8730 12469 8732
rect 12493 8730 12549 8732
rect 12253 8678 12299 8730
rect 12299 8678 12309 8730
rect 12333 8678 12363 8730
rect 12363 8678 12375 8730
rect 12375 8678 12389 8730
rect 12413 8678 12427 8730
rect 12427 8678 12439 8730
rect 12439 8678 12469 8730
rect 12493 8678 12503 8730
rect 12503 8678 12549 8730
rect 12253 8676 12309 8678
rect 12333 8676 12389 8678
rect 12413 8676 12469 8678
rect 12493 8676 12549 8678
rect 12530 7828 12532 7848
rect 12532 7828 12584 7848
rect 12584 7828 12586 7848
rect 12530 7792 12586 7828
rect 12253 7642 12309 7644
rect 12333 7642 12389 7644
rect 12413 7642 12469 7644
rect 12493 7642 12549 7644
rect 12253 7590 12299 7642
rect 12299 7590 12309 7642
rect 12333 7590 12363 7642
rect 12363 7590 12375 7642
rect 12375 7590 12389 7642
rect 12413 7590 12427 7642
rect 12427 7590 12439 7642
rect 12439 7590 12469 7642
rect 12493 7590 12503 7642
rect 12503 7590 12549 7642
rect 12253 7588 12309 7590
rect 12333 7588 12389 7590
rect 12413 7588 12469 7590
rect 12493 7588 12549 7590
rect 11978 7404 12034 7440
rect 11978 7384 11980 7404
rect 11980 7384 12032 7404
rect 12032 7384 12034 7404
rect 11593 7098 11649 7100
rect 11673 7098 11729 7100
rect 11753 7098 11809 7100
rect 11833 7098 11889 7100
rect 11593 7046 11639 7098
rect 11639 7046 11649 7098
rect 11673 7046 11703 7098
rect 11703 7046 11715 7098
rect 11715 7046 11729 7098
rect 11753 7046 11767 7098
rect 11767 7046 11779 7098
rect 11779 7046 11809 7098
rect 11833 7046 11843 7098
rect 11843 7046 11889 7098
rect 11593 7044 11649 7046
rect 11673 7044 11729 7046
rect 11753 7044 11809 7046
rect 11833 7044 11889 7046
rect 11886 6740 11888 6760
rect 11888 6740 11940 6760
rect 11940 6740 11942 6760
rect 11886 6704 11942 6740
rect 11886 6296 11942 6352
rect 11242 5652 11244 5672
rect 11244 5652 11296 5672
rect 11296 5652 11298 5672
rect 11242 5616 11298 5652
rect 11593 6010 11649 6012
rect 11673 6010 11729 6012
rect 11753 6010 11809 6012
rect 11833 6010 11889 6012
rect 11593 5958 11639 6010
rect 11639 5958 11649 6010
rect 11673 5958 11703 6010
rect 11703 5958 11715 6010
rect 11715 5958 11729 6010
rect 11753 5958 11767 6010
rect 11767 5958 11779 6010
rect 11779 5958 11809 6010
rect 11833 5958 11843 6010
rect 11843 5958 11889 6010
rect 11593 5956 11649 5958
rect 11673 5956 11729 5958
rect 11753 5956 11809 5958
rect 11833 5956 11889 5958
rect 11593 4922 11649 4924
rect 11673 4922 11729 4924
rect 11753 4922 11809 4924
rect 11833 4922 11889 4924
rect 11593 4870 11639 4922
rect 11639 4870 11649 4922
rect 11673 4870 11703 4922
rect 11703 4870 11715 4922
rect 11715 4870 11729 4922
rect 11753 4870 11767 4922
rect 11767 4870 11779 4922
rect 11779 4870 11809 4922
rect 11833 4870 11843 4922
rect 11843 4870 11889 4922
rect 11593 4868 11649 4870
rect 11673 4868 11729 4870
rect 11753 4868 11809 4870
rect 11833 4868 11889 4870
rect 11593 3834 11649 3836
rect 11673 3834 11729 3836
rect 11753 3834 11809 3836
rect 11833 3834 11889 3836
rect 11593 3782 11639 3834
rect 11639 3782 11649 3834
rect 11673 3782 11703 3834
rect 11703 3782 11715 3834
rect 11715 3782 11729 3834
rect 11753 3782 11767 3834
rect 11767 3782 11779 3834
rect 11779 3782 11809 3834
rect 11833 3782 11843 3834
rect 11843 3782 11889 3834
rect 11593 3780 11649 3782
rect 11673 3780 11729 3782
rect 11753 3780 11809 3782
rect 11833 3780 11889 3782
rect 11593 2746 11649 2748
rect 11673 2746 11729 2748
rect 11753 2746 11809 2748
rect 11833 2746 11889 2748
rect 11593 2694 11639 2746
rect 11639 2694 11649 2746
rect 11673 2694 11703 2746
rect 11703 2694 11715 2746
rect 11715 2694 11729 2746
rect 11753 2694 11767 2746
rect 11767 2694 11779 2746
rect 11779 2694 11809 2746
rect 11833 2694 11843 2746
rect 11843 2694 11889 2746
rect 11593 2692 11649 2694
rect 11673 2692 11729 2694
rect 11753 2692 11809 2694
rect 11833 2692 11889 2694
rect 12806 10260 12862 10296
rect 12806 10240 12808 10260
rect 12808 10240 12860 10260
rect 12860 10240 12862 10260
rect 13818 14728 13874 14784
rect 16508 18522 16564 18524
rect 16588 18522 16644 18524
rect 16668 18522 16724 18524
rect 16748 18522 16804 18524
rect 16508 18470 16554 18522
rect 16554 18470 16564 18522
rect 16588 18470 16618 18522
rect 16618 18470 16630 18522
rect 16630 18470 16644 18522
rect 16668 18470 16682 18522
rect 16682 18470 16694 18522
rect 16694 18470 16724 18522
rect 16748 18470 16758 18522
rect 16758 18470 16804 18522
rect 16508 18468 16564 18470
rect 16588 18468 16644 18470
rect 16668 18468 16724 18470
rect 16748 18468 16804 18470
rect 14370 14728 14426 14784
rect 15848 17978 15904 17980
rect 15928 17978 15984 17980
rect 16008 17978 16064 17980
rect 16088 17978 16144 17980
rect 15848 17926 15894 17978
rect 15894 17926 15904 17978
rect 15928 17926 15958 17978
rect 15958 17926 15970 17978
rect 15970 17926 15984 17978
rect 16008 17926 16022 17978
rect 16022 17926 16034 17978
rect 16034 17926 16064 17978
rect 16088 17926 16098 17978
rect 16098 17926 16144 17978
rect 15848 17924 15904 17926
rect 15928 17924 15984 17926
rect 16008 17924 16064 17926
rect 16088 17924 16144 17926
rect 15848 16890 15904 16892
rect 15928 16890 15984 16892
rect 16008 16890 16064 16892
rect 16088 16890 16144 16892
rect 15848 16838 15894 16890
rect 15894 16838 15904 16890
rect 15928 16838 15958 16890
rect 15958 16838 15970 16890
rect 15970 16838 15984 16890
rect 16008 16838 16022 16890
rect 16022 16838 16034 16890
rect 16034 16838 16064 16890
rect 16088 16838 16098 16890
rect 16098 16838 16144 16890
rect 15848 16836 15904 16838
rect 15928 16836 15984 16838
rect 16008 16836 16064 16838
rect 16088 16836 16144 16838
rect 13726 13776 13782 13832
rect 13358 10004 13360 10024
rect 13360 10004 13412 10024
rect 13412 10004 13414 10024
rect 13358 9968 13414 10004
rect 12253 6554 12309 6556
rect 12333 6554 12389 6556
rect 12413 6554 12469 6556
rect 12493 6554 12549 6556
rect 12253 6502 12299 6554
rect 12299 6502 12309 6554
rect 12333 6502 12363 6554
rect 12363 6502 12375 6554
rect 12375 6502 12389 6554
rect 12413 6502 12427 6554
rect 12427 6502 12439 6554
rect 12439 6502 12469 6554
rect 12493 6502 12503 6554
rect 12503 6502 12549 6554
rect 12253 6500 12309 6502
rect 12333 6500 12389 6502
rect 12413 6500 12469 6502
rect 12493 6500 12549 6502
rect 12253 5466 12309 5468
rect 12333 5466 12389 5468
rect 12413 5466 12469 5468
rect 12493 5466 12549 5468
rect 12253 5414 12299 5466
rect 12299 5414 12309 5466
rect 12333 5414 12363 5466
rect 12363 5414 12375 5466
rect 12375 5414 12389 5466
rect 12413 5414 12427 5466
rect 12427 5414 12439 5466
rect 12439 5414 12469 5466
rect 12493 5414 12503 5466
rect 12503 5414 12549 5466
rect 12253 5412 12309 5414
rect 12333 5412 12389 5414
rect 12413 5412 12469 5414
rect 12493 5412 12549 5414
rect 12253 4378 12309 4380
rect 12333 4378 12389 4380
rect 12413 4378 12469 4380
rect 12493 4378 12549 4380
rect 12253 4326 12299 4378
rect 12299 4326 12309 4378
rect 12333 4326 12363 4378
rect 12363 4326 12375 4378
rect 12375 4326 12389 4378
rect 12413 4326 12427 4378
rect 12427 4326 12439 4378
rect 12439 4326 12469 4378
rect 12493 4326 12503 4378
rect 12503 4326 12549 4378
rect 12253 4324 12309 4326
rect 12333 4324 12389 4326
rect 12413 4324 12469 4326
rect 12493 4324 12549 4326
rect 12253 3290 12309 3292
rect 12333 3290 12389 3292
rect 12413 3290 12469 3292
rect 12493 3290 12549 3292
rect 12253 3238 12299 3290
rect 12299 3238 12309 3290
rect 12333 3238 12363 3290
rect 12363 3238 12375 3290
rect 12375 3238 12389 3290
rect 12413 3238 12427 3290
rect 12427 3238 12439 3290
rect 12439 3238 12469 3290
rect 12493 3238 12503 3290
rect 12503 3238 12549 3290
rect 12253 3236 12309 3238
rect 12333 3236 12389 3238
rect 12413 3236 12469 3238
rect 12493 3236 12549 3238
rect 13910 9968 13966 10024
rect 15848 15802 15904 15804
rect 15928 15802 15984 15804
rect 16008 15802 16064 15804
rect 16088 15802 16144 15804
rect 15848 15750 15894 15802
rect 15894 15750 15904 15802
rect 15928 15750 15958 15802
rect 15958 15750 15970 15802
rect 15970 15750 15984 15802
rect 16008 15750 16022 15802
rect 16022 15750 16034 15802
rect 16034 15750 16064 15802
rect 16088 15750 16098 15802
rect 16098 15750 16144 15802
rect 15848 15748 15904 15750
rect 15928 15748 15984 15750
rect 16008 15748 16064 15750
rect 16088 15748 16144 15750
rect 16508 17434 16564 17436
rect 16588 17434 16644 17436
rect 16668 17434 16724 17436
rect 16748 17434 16804 17436
rect 16508 17382 16554 17434
rect 16554 17382 16564 17434
rect 16588 17382 16618 17434
rect 16618 17382 16630 17434
rect 16630 17382 16644 17434
rect 16668 17382 16682 17434
rect 16682 17382 16694 17434
rect 16694 17382 16724 17434
rect 16748 17382 16758 17434
rect 16758 17382 16804 17434
rect 16508 17380 16564 17382
rect 16588 17380 16644 17382
rect 16668 17380 16724 17382
rect 16748 17380 16804 17382
rect 16508 16346 16564 16348
rect 16588 16346 16644 16348
rect 16668 16346 16724 16348
rect 16748 16346 16804 16348
rect 16508 16294 16554 16346
rect 16554 16294 16564 16346
rect 16588 16294 16618 16346
rect 16618 16294 16630 16346
rect 16630 16294 16644 16346
rect 16668 16294 16682 16346
rect 16682 16294 16694 16346
rect 16694 16294 16724 16346
rect 16748 16294 16758 16346
rect 16758 16294 16804 16346
rect 16508 16292 16564 16294
rect 16588 16292 16644 16294
rect 16668 16292 16724 16294
rect 16748 16292 16804 16294
rect 17682 15680 17738 15736
rect 16508 15258 16564 15260
rect 16588 15258 16644 15260
rect 16668 15258 16724 15260
rect 16748 15258 16804 15260
rect 16508 15206 16554 15258
rect 16554 15206 16564 15258
rect 16588 15206 16618 15258
rect 16618 15206 16630 15258
rect 16630 15206 16644 15258
rect 16668 15206 16682 15258
rect 16682 15206 16694 15258
rect 16694 15206 16724 15258
rect 16748 15206 16758 15258
rect 16758 15206 16804 15258
rect 16508 15204 16564 15206
rect 16588 15204 16644 15206
rect 16668 15204 16724 15206
rect 16748 15204 16804 15206
rect 15848 14714 15904 14716
rect 15928 14714 15984 14716
rect 16008 14714 16064 14716
rect 16088 14714 16144 14716
rect 15848 14662 15894 14714
rect 15894 14662 15904 14714
rect 15928 14662 15958 14714
rect 15958 14662 15970 14714
rect 15970 14662 15984 14714
rect 16008 14662 16022 14714
rect 16022 14662 16034 14714
rect 16034 14662 16064 14714
rect 16088 14662 16098 14714
rect 16098 14662 16144 14714
rect 15848 14660 15904 14662
rect 15928 14660 15984 14662
rect 16008 14660 16064 14662
rect 16088 14660 16144 14662
rect 14370 7928 14426 7984
rect 14002 6296 14058 6352
rect 14554 7792 14610 7848
rect 14370 5772 14426 5808
rect 14370 5752 14372 5772
rect 14372 5752 14424 5772
rect 14424 5752 14426 5772
rect 15848 13626 15904 13628
rect 15928 13626 15984 13628
rect 16008 13626 16064 13628
rect 16088 13626 16144 13628
rect 15848 13574 15894 13626
rect 15894 13574 15904 13626
rect 15928 13574 15958 13626
rect 15958 13574 15970 13626
rect 15970 13574 15984 13626
rect 16008 13574 16022 13626
rect 16022 13574 16034 13626
rect 16034 13574 16064 13626
rect 16088 13574 16098 13626
rect 16098 13574 16144 13626
rect 15848 13572 15904 13574
rect 15928 13572 15984 13574
rect 16008 13572 16064 13574
rect 16088 13572 16144 13574
rect 16946 14320 17002 14376
rect 16508 14170 16564 14172
rect 16588 14170 16644 14172
rect 16668 14170 16724 14172
rect 16748 14170 16804 14172
rect 16508 14118 16554 14170
rect 16554 14118 16564 14170
rect 16588 14118 16618 14170
rect 16618 14118 16630 14170
rect 16630 14118 16644 14170
rect 16668 14118 16682 14170
rect 16682 14118 16694 14170
rect 16694 14118 16724 14170
rect 16748 14118 16758 14170
rect 16758 14118 16804 14170
rect 16508 14116 16564 14118
rect 16588 14116 16644 14118
rect 16668 14116 16724 14118
rect 16748 14116 16804 14118
rect 15848 12538 15904 12540
rect 15928 12538 15984 12540
rect 16008 12538 16064 12540
rect 16088 12538 16144 12540
rect 15848 12486 15894 12538
rect 15894 12486 15904 12538
rect 15928 12486 15958 12538
rect 15958 12486 15970 12538
rect 15970 12486 15984 12538
rect 16008 12486 16022 12538
rect 16022 12486 16034 12538
rect 16034 12486 16064 12538
rect 16088 12486 16098 12538
rect 16098 12486 16144 12538
rect 15848 12484 15904 12486
rect 15928 12484 15984 12486
rect 16008 12484 16064 12486
rect 16088 12484 16144 12486
rect 17682 15000 17738 15056
rect 16508 13082 16564 13084
rect 16588 13082 16644 13084
rect 16668 13082 16724 13084
rect 16748 13082 16804 13084
rect 16508 13030 16554 13082
rect 16554 13030 16564 13082
rect 16588 13030 16618 13082
rect 16618 13030 16630 13082
rect 16630 13030 16644 13082
rect 16668 13030 16682 13082
rect 16682 13030 16694 13082
rect 16694 13030 16724 13082
rect 16748 13030 16758 13082
rect 16758 13030 16804 13082
rect 16508 13028 16564 13030
rect 16588 13028 16644 13030
rect 16668 13028 16724 13030
rect 16748 13028 16804 13030
rect 16302 12436 16358 12472
rect 16302 12416 16304 12436
rect 16304 12416 16356 12436
rect 16356 12416 16358 12436
rect 16578 12416 16634 12472
rect 15848 11450 15904 11452
rect 15928 11450 15984 11452
rect 16008 11450 16064 11452
rect 16088 11450 16144 11452
rect 15848 11398 15894 11450
rect 15894 11398 15904 11450
rect 15928 11398 15958 11450
rect 15958 11398 15970 11450
rect 15970 11398 15984 11450
rect 16008 11398 16022 11450
rect 16022 11398 16034 11450
rect 16034 11398 16064 11450
rect 16088 11398 16098 11450
rect 16098 11398 16144 11450
rect 15848 11396 15904 11398
rect 15928 11396 15984 11398
rect 16008 11396 16064 11398
rect 16088 11396 16144 11398
rect 16508 11994 16564 11996
rect 16588 11994 16644 11996
rect 16668 11994 16724 11996
rect 16748 11994 16804 11996
rect 16508 11942 16554 11994
rect 16554 11942 16564 11994
rect 16588 11942 16618 11994
rect 16618 11942 16630 11994
rect 16630 11942 16644 11994
rect 16668 11942 16682 11994
rect 16682 11942 16694 11994
rect 16694 11942 16724 11994
rect 16748 11942 16758 11994
rect 16758 11942 16804 11994
rect 16508 11940 16564 11942
rect 16588 11940 16644 11942
rect 16668 11940 16724 11942
rect 16748 11940 16804 11942
rect 16508 10906 16564 10908
rect 16588 10906 16644 10908
rect 16668 10906 16724 10908
rect 16748 10906 16804 10908
rect 16508 10854 16554 10906
rect 16554 10854 16564 10906
rect 16588 10854 16618 10906
rect 16618 10854 16630 10906
rect 16630 10854 16644 10906
rect 16668 10854 16682 10906
rect 16682 10854 16694 10906
rect 16694 10854 16724 10906
rect 16748 10854 16758 10906
rect 16758 10854 16804 10906
rect 16508 10852 16564 10854
rect 16588 10852 16644 10854
rect 16668 10852 16724 10854
rect 16748 10852 16804 10854
rect 15848 10362 15904 10364
rect 15928 10362 15984 10364
rect 16008 10362 16064 10364
rect 16088 10362 16144 10364
rect 15848 10310 15894 10362
rect 15894 10310 15904 10362
rect 15928 10310 15958 10362
rect 15958 10310 15970 10362
rect 15970 10310 15984 10362
rect 16008 10310 16022 10362
rect 16022 10310 16034 10362
rect 16034 10310 16064 10362
rect 16088 10310 16098 10362
rect 16098 10310 16144 10362
rect 15848 10308 15904 10310
rect 15928 10308 15984 10310
rect 16008 10308 16064 10310
rect 16088 10308 16144 10310
rect 15014 9968 15070 10024
rect 16508 9818 16564 9820
rect 16588 9818 16644 9820
rect 16668 9818 16724 9820
rect 16748 9818 16804 9820
rect 16508 9766 16554 9818
rect 16554 9766 16564 9818
rect 16588 9766 16618 9818
rect 16618 9766 16630 9818
rect 16630 9766 16644 9818
rect 16668 9766 16682 9818
rect 16682 9766 16694 9818
rect 16694 9766 16724 9818
rect 16748 9766 16758 9818
rect 16758 9766 16804 9818
rect 16508 9764 16564 9766
rect 16588 9764 16644 9766
rect 16668 9764 16724 9766
rect 16748 9764 16804 9766
rect 14922 7384 14978 7440
rect 14462 5616 14518 5672
rect 14830 6840 14886 6896
rect 15848 9274 15904 9276
rect 15928 9274 15984 9276
rect 16008 9274 16064 9276
rect 16088 9274 16144 9276
rect 15848 9222 15894 9274
rect 15894 9222 15904 9274
rect 15928 9222 15958 9274
rect 15958 9222 15970 9274
rect 15970 9222 15984 9274
rect 16008 9222 16022 9274
rect 16022 9222 16034 9274
rect 16034 9222 16064 9274
rect 16088 9222 16098 9274
rect 16098 9222 16144 9274
rect 15848 9220 15904 9222
rect 15928 9220 15984 9222
rect 16008 9220 16064 9222
rect 16088 9220 16144 9222
rect 15848 8186 15904 8188
rect 15928 8186 15984 8188
rect 16008 8186 16064 8188
rect 16088 8186 16144 8188
rect 15848 8134 15894 8186
rect 15894 8134 15904 8186
rect 15928 8134 15958 8186
rect 15958 8134 15970 8186
rect 15970 8134 15984 8186
rect 16008 8134 16022 8186
rect 16022 8134 16034 8186
rect 16034 8134 16064 8186
rect 16088 8134 16098 8186
rect 16098 8134 16144 8186
rect 15848 8132 15904 8134
rect 15928 8132 15984 8134
rect 16008 8132 16064 8134
rect 16088 8132 16144 8134
rect 15848 7098 15904 7100
rect 15928 7098 15984 7100
rect 16008 7098 16064 7100
rect 16088 7098 16144 7100
rect 15848 7046 15894 7098
rect 15894 7046 15904 7098
rect 15928 7046 15958 7098
rect 15958 7046 15970 7098
rect 15970 7046 15984 7098
rect 16008 7046 16022 7098
rect 16022 7046 16034 7098
rect 16034 7046 16064 7098
rect 16088 7046 16098 7098
rect 16098 7046 16144 7098
rect 15848 7044 15904 7046
rect 15928 7044 15984 7046
rect 16008 7044 16064 7046
rect 16088 7044 16144 7046
rect 17682 12960 17738 13016
rect 16508 8730 16564 8732
rect 16588 8730 16644 8732
rect 16668 8730 16724 8732
rect 16748 8730 16804 8732
rect 16508 8678 16554 8730
rect 16554 8678 16564 8730
rect 16588 8678 16618 8730
rect 16618 8678 16630 8730
rect 16630 8678 16644 8730
rect 16668 8678 16682 8730
rect 16682 8678 16694 8730
rect 16694 8678 16724 8730
rect 16748 8678 16758 8730
rect 16758 8678 16804 8730
rect 16508 8676 16564 8678
rect 16588 8676 16644 8678
rect 16668 8676 16724 8678
rect 16748 8676 16804 8678
rect 17682 10240 17738 10296
rect 16946 8200 17002 8256
rect 16508 7642 16564 7644
rect 16588 7642 16644 7644
rect 16668 7642 16724 7644
rect 16748 7642 16804 7644
rect 16508 7590 16554 7642
rect 16554 7590 16564 7642
rect 16588 7590 16618 7642
rect 16618 7590 16630 7642
rect 16630 7590 16644 7642
rect 16668 7590 16682 7642
rect 16682 7590 16694 7642
rect 16694 7590 16724 7642
rect 16748 7590 16758 7642
rect 16758 7590 16804 7642
rect 16508 7588 16564 7590
rect 16588 7588 16644 7590
rect 16668 7588 16724 7590
rect 16748 7588 16804 7590
rect 17774 7520 17830 7576
rect 17774 6840 17830 6896
rect 15848 6010 15904 6012
rect 15928 6010 15984 6012
rect 16008 6010 16064 6012
rect 16088 6010 16144 6012
rect 15848 5958 15894 6010
rect 15894 5958 15904 6010
rect 15928 5958 15958 6010
rect 15958 5958 15970 6010
rect 15970 5958 15984 6010
rect 16008 5958 16022 6010
rect 16022 5958 16034 6010
rect 16034 5958 16064 6010
rect 16088 5958 16098 6010
rect 16098 5958 16144 6010
rect 15848 5956 15904 5958
rect 15928 5956 15984 5958
rect 16008 5956 16064 5958
rect 16088 5956 16144 5958
rect 15848 4922 15904 4924
rect 15928 4922 15984 4924
rect 16008 4922 16064 4924
rect 16088 4922 16144 4924
rect 15848 4870 15894 4922
rect 15894 4870 15904 4922
rect 15928 4870 15958 4922
rect 15958 4870 15970 4922
rect 15970 4870 15984 4922
rect 16008 4870 16022 4922
rect 16022 4870 16034 4922
rect 16034 4870 16064 4922
rect 16088 4870 16098 4922
rect 16098 4870 16144 4922
rect 15848 4868 15904 4870
rect 15928 4868 15984 4870
rect 16008 4868 16064 4870
rect 16088 4868 16144 4870
rect 16508 6554 16564 6556
rect 16588 6554 16644 6556
rect 16668 6554 16724 6556
rect 16748 6554 16804 6556
rect 16508 6502 16554 6554
rect 16554 6502 16564 6554
rect 16588 6502 16618 6554
rect 16618 6502 16630 6554
rect 16630 6502 16644 6554
rect 16668 6502 16682 6554
rect 16682 6502 16694 6554
rect 16694 6502 16724 6554
rect 16748 6502 16758 6554
rect 16758 6502 16804 6554
rect 16508 6500 16564 6502
rect 16588 6500 16644 6502
rect 16668 6500 16724 6502
rect 16748 6500 16804 6502
rect 16508 5466 16564 5468
rect 16588 5466 16644 5468
rect 16668 5466 16724 5468
rect 16748 5466 16804 5468
rect 16508 5414 16554 5466
rect 16554 5414 16564 5466
rect 16588 5414 16618 5466
rect 16618 5414 16630 5466
rect 16630 5414 16644 5466
rect 16668 5414 16682 5466
rect 16682 5414 16694 5466
rect 16694 5414 16724 5466
rect 16748 5414 16758 5466
rect 16758 5414 16804 5466
rect 16508 5412 16564 5414
rect 16588 5412 16644 5414
rect 16668 5412 16724 5414
rect 16748 5412 16804 5414
rect 16508 4378 16564 4380
rect 16588 4378 16644 4380
rect 16668 4378 16724 4380
rect 16748 4378 16804 4380
rect 16508 4326 16554 4378
rect 16554 4326 16564 4378
rect 16588 4326 16618 4378
rect 16618 4326 16630 4378
rect 16630 4326 16644 4378
rect 16668 4326 16682 4378
rect 16682 4326 16694 4378
rect 16694 4326 16724 4378
rect 16748 4326 16758 4378
rect 16758 4326 16804 4378
rect 16508 4324 16564 4326
rect 16588 4324 16644 4326
rect 16668 4324 16724 4326
rect 16748 4324 16804 4326
rect 17774 6160 17830 6216
rect 17682 5480 17738 5536
rect 17590 4800 17646 4856
rect 15848 3834 15904 3836
rect 15928 3834 15984 3836
rect 16008 3834 16064 3836
rect 16088 3834 16144 3836
rect 15848 3782 15894 3834
rect 15894 3782 15904 3834
rect 15928 3782 15958 3834
rect 15958 3782 15970 3834
rect 15970 3782 15984 3834
rect 16008 3782 16022 3834
rect 16022 3782 16034 3834
rect 16034 3782 16064 3834
rect 16088 3782 16098 3834
rect 16098 3782 16144 3834
rect 15848 3780 15904 3782
rect 15928 3780 15984 3782
rect 16008 3780 16064 3782
rect 16088 3780 16144 3782
rect 14646 2896 14702 2952
rect 17682 3460 17738 3496
rect 17682 3440 17684 3460
rect 17684 3440 17736 3460
rect 17736 3440 17738 3460
rect 16508 3290 16564 3292
rect 16588 3290 16644 3292
rect 16668 3290 16724 3292
rect 16748 3290 16804 3292
rect 16508 3238 16554 3290
rect 16554 3238 16564 3290
rect 16588 3238 16618 3290
rect 16618 3238 16630 3290
rect 16630 3238 16644 3290
rect 16668 3238 16682 3290
rect 16682 3238 16694 3290
rect 16694 3238 16724 3290
rect 16748 3238 16758 3290
rect 16758 3238 16804 3290
rect 16508 3236 16564 3238
rect 16588 3236 16644 3238
rect 16668 3236 16724 3238
rect 16748 3236 16804 3238
rect 15848 2746 15904 2748
rect 15928 2746 15984 2748
rect 16008 2746 16064 2748
rect 16088 2746 16144 2748
rect 15848 2694 15894 2746
rect 15894 2694 15904 2746
rect 15928 2694 15958 2746
rect 15958 2694 15970 2746
rect 15970 2694 15984 2746
rect 16008 2694 16022 2746
rect 16022 2694 16034 2746
rect 16034 2694 16064 2746
rect 16088 2694 16098 2746
rect 16098 2694 16144 2746
rect 15848 2692 15904 2694
rect 15928 2692 15984 2694
rect 16008 2692 16064 2694
rect 16088 2692 16144 2694
rect 12253 2202 12309 2204
rect 12333 2202 12389 2204
rect 12413 2202 12469 2204
rect 12493 2202 12549 2204
rect 12253 2150 12299 2202
rect 12299 2150 12309 2202
rect 12333 2150 12363 2202
rect 12363 2150 12375 2202
rect 12375 2150 12389 2202
rect 12413 2150 12427 2202
rect 12427 2150 12439 2202
rect 12439 2150 12469 2202
rect 12493 2150 12503 2202
rect 12503 2150 12549 2202
rect 12253 2148 12309 2150
rect 12333 2148 12389 2150
rect 12413 2148 12469 2150
rect 12493 2148 12549 2150
rect 16508 2202 16564 2204
rect 16588 2202 16644 2204
rect 16668 2202 16724 2204
rect 16748 2202 16804 2204
rect 16508 2150 16554 2202
rect 16554 2150 16564 2202
rect 16588 2150 16618 2202
rect 16618 2150 16630 2202
rect 16630 2150 16644 2202
rect 16668 2150 16682 2202
rect 16682 2150 16694 2202
rect 16694 2150 16724 2202
rect 16748 2150 16758 2202
rect 16758 2150 16804 2202
rect 16508 2148 16564 2150
rect 16588 2148 16644 2150
rect 16668 2148 16724 2150
rect 16748 2148 16804 2150
<< metal3 >>
rect 3073 19072 3389 19073
rect 3073 19008 3079 19072
rect 3143 19008 3159 19072
rect 3223 19008 3239 19072
rect 3303 19008 3319 19072
rect 3383 19008 3389 19072
rect 3073 19007 3389 19008
rect 7328 19072 7644 19073
rect 7328 19008 7334 19072
rect 7398 19008 7414 19072
rect 7478 19008 7494 19072
rect 7558 19008 7574 19072
rect 7638 19008 7644 19072
rect 7328 19007 7644 19008
rect 11583 19072 11899 19073
rect 11583 19008 11589 19072
rect 11653 19008 11669 19072
rect 11733 19008 11749 19072
rect 11813 19008 11829 19072
rect 11893 19008 11899 19072
rect 11583 19007 11899 19008
rect 15838 19072 16154 19073
rect 15838 19008 15844 19072
rect 15908 19008 15924 19072
rect 15988 19008 16004 19072
rect 16068 19008 16084 19072
rect 16148 19008 16154 19072
rect 15838 19007 16154 19008
rect 3733 18528 4049 18529
rect 3733 18464 3739 18528
rect 3803 18464 3819 18528
rect 3883 18464 3899 18528
rect 3963 18464 3979 18528
rect 4043 18464 4049 18528
rect 3733 18463 4049 18464
rect 7988 18528 8304 18529
rect 7988 18464 7994 18528
rect 8058 18464 8074 18528
rect 8138 18464 8154 18528
rect 8218 18464 8234 18528
rect 8298 18464 8304 18528
rect 7988 18463 8304 18464
rect 12243 18528 12559 18529
rect 12243 18464 12249 18528
rect 12313 18464 12329 18528
rect 12393 18464 12409 18528
rect 12473 18464 12489 18528
rect 12553 18464 12559 18528
rect 12243 18463 12559 18464
rect 16498 18528 16814 18529
rect 16498 18464 16504 18528
rect 16568 18464 16584 18528
rect 16648 18464 16664 18528
rect 16728 18464 16744 18528
rect 16808 18464 16814 18528
rect 16498 18463 16814 18464
rect 3073 17984 3389 17985
rect 3073 17920 3079 17984
rect 3143 17920 3159 17984
rect 3223 17920 3239 17984
rect 3303 17920 3319 17984
rect 3383 17920 3389 17984
rect 3073 17919 3389 17920
rect 7328 17984 7644 17985
rect 7328 17920 7334 17984
rect 7398 17920 7414 17984
rect 7478 17920 7494 17984
rect 7558 17920 7574 17984
rect 7638 17920 7644 17984
rect 7328 17919 7644 17920
rect 11583 17984 11899 17985
rect 11583 17920 11589 17984
rect 11653 17920 11669 17984
rect 11733 17920 11749 17984
rect 11813 17920 11829 17984
rect 11893 17920 11899 17984
rect 11583 17919 11899 17920
rect 15838 17984 16154 17985
rect 15838 17920 15844 17984
rect 15908 17920 15924 17984
rect 15988 17920 16004 17984
rect 16068 17920 16084 17984
rect 16148 17920 16154 17984
rect 15838 17919 16154 17920
rect 0 17778 800 17808
rect 3550 17778 3556 17780
rect 0 17718 3556 17778
rect 0 17688 800 17718
rect 3550 17716 3556 17718
rect 3620 17716 3626 17780
rect 3733 17440 4049 17441
rect 3733 17376 3739 17440
rect 3803 17376 3819 17440
rect 3883 17376 3899 17440
rect 3963 17376 3979 17440
rect 4043 17376 4049 17440
rect 3733 17375 4049 17376
rect 7988 17440 8304 17441
rect 7988 17376 7994 17440
rect 8058 17376 8074 17440
rect 8138 17376 8154 17440
rect 8218 17376 8234 17440
rect 8298 17376 8304 17440
rect 7988 17375 8304 17376
rect 12243 17440 12559 17441
rect 12243 17376 12249 17440
rect 12313 17376 12329 17440
rect 12393 17376 12409 17440
rect 12473 17376 12489 17440
rect 12553 17376 12559 17440
rect 12243 17375 12559 17376
rect 16498 17440 16814 17441
rect 16498 17376 16504 17440
rect 16568 17376 16584 17440
rect 16648 17376 16664 17440
rect 16728 17376 16744 17440
rect 16808 17376 16814 17440
rect 16498 17375 16814 17376
rect 3073 16896 3389 16897
rect 3073 16832 3079 16896
rect 3143 16832 3159 16896
rect 3223 16832 3239 16896
rect 3303 16832 3319 16896
rect 3383 16832 3389 16896
rect 3073 16831 3389 16832
rect 7328 16896 7644 16897
rect 7328 16832 7334 16896
rect 7398 16832 7414 16896
rect 7478 16832 7494 16896
rect 7558 16832 7574 16896
rect 7638 16832 7644 16896
rect 7328 16831 7644 16832
rect 11583 16896 11899 16897
rect 11583 16832 11589 16896
rect 11653 16832 11669 16896
rect 11733 16832 11749 16896
rect 11813 16832 11829 16896
rect 11893 16832 11899 16896
rect 11583 16831 11899 16832
rect 15838 16896 16154 16897
rect 15838 16832 15844 16896
rect 15908 16832 15924 16896
rect 15988 16832 16004 16896
rect 16068 16832 16084 16896
rect 16148 16832 16154 16896
rect 15838 16831 16154 16832
rect 841 16554 907 16557
rect 798 16552 907 16554
rect 798 16496 846 16552
rect 902 16496 907 16552
rect 798 16491 907 16496
rect 798 16448 858 16491
rect 0 16358 858 16448
rect 0 16328 800 16358
rect 3733 16352 4049 16353
rect 3733 16288 3739 16352
rect 3803 16288 3819 16352
rect 3883 16288 3899 16352
rect 3963 16288 3979 16352
rect 4043 16288 4049 16352
rect 3733 16287 4049 16288
rect 7988 16352 8304 16353
rect 7988 16288 7994 16352
rect 8058 16288 8074 16352
rect 8138 16288 8154 16352
rect 8218 16288 8234 16352
rect 8298 16288 8304 16352
rect 7988 16287 8304 16288
rect 12243 16352 12559 16353
rect 12243 16288 12249 16352
rect 12313 16288 12329 16352
rect 12393 16288 12409 16352
rect 12473 16288 12489 16352
rect 12553 16288 12559 16352
rect 12243 16287 12559 16288
rect 16498 16352 16814 16353
rect 16498 16288 16504 16352
rect 16568 16288 16584 16352
rect 16648 16288 16664 16352
rect 16728 16288 16744 16352
rect 16808 16288 16814 16352
rect 16498 16287 16814 16288
rect 3073 15808 3389 15809
rect 3073 15744 3079 15808
rect 3143 15744 3159 15808
rect 3223 15744 3239 15808
rect 3303 15744 3319 15808
rect 3383 15744 3389 15808
rect 3073 15743 3389 15744
rect 7328 15808 7644 15809
rect 7328 15744 7334 15808
rect 7398 15744 7414 15808
rect 7478 15744 7494 15808
rect 7558 15744 7574 15808
rect 7638 15744 7644 15808
rect 7328 15743 7644 15744
rect 11583 15808 11899 15809
rect 11583 15744 11589 15808
rect 11653 15744 11669 15808
rect 11733 15744 11749 15808
rect 11813 15744 11829 15808
rect 11893 15744 11899 15808
rect 11583 15743 11899 15744
rect 15838 15808 16154 15809
rect 15838 15744 15844 15808
rect 15908 15744 15924 15808
rect 15988 15744 16004 15808
rect 16068 15744 16084 15808
rect 16148 15744 16154 15808
rect 15838 15743 16154 15744
rect 17677 15738 17743 15741
rect 18469 15738 19269 15768
rect 17677 15736 19269 15738
rect 17677 15680 17682 15736
rect 17738 15680 19269 15736
rect 17677 15678 19269 15680
rect 17677 15675 17743 15678
rect 18469 15648 19269 15678
rect 3733 15264 4049 15265
rect 3733 15200 3739 15264
rect 3803 15200 3819 15264
rect 3883 15200 3899 15264
rect 3963 15200 3979 15264
rect 4043 15200 4049 15264
rect 3733 15199 4049 15200
rect 7988 15264 8304 15265
rect 7988 15200 7994 15264
rect 8058 15200 8074 15264
rect 8138 15200 8154 15264
rect 8218 15200 8234 15264
rect 8298 15200 8304 15264
rect 7988 15199 8304 15200
rect 12243 15264 12559 15265
rect 12243 15200 12249 15264
rect 12313 15200 12329 15264
rect 12393 15200 12409 15264
rect 12473 15200 12489 15264
rect 12553 15200 12559 15264
rect 12243 15199 12559 15200
rect 16498 15264 16814 15265
rect 16498 15200 16504 15264
rect 16568 15200 16584 15264
rect 16648 15200 16664 15264
rect 16728 15200 16744 15264
rect 16808 15200 16814 15264
rect 16498 15199 16814 15200
rect 0 15058 800 15088
rect 1485 15058 1551 15061
rect 12709 15060 12775 15061
rect 12709 15058 12756 15060
rect 0 15056 1551 15058
rect 0 15000 1490 15056
rect 1546 15000 1551 15056
rect 0 14998 1551 15000
rect 12664 15056 12756 15058
rect 12664 15000 12714 15056
rect 12664 14998 12756 15000
rect 0 14968 800 14998
rect 1485 14995 1551 14998
rect 12709 14996 12756 14998
rect 12820 14996 12826 15060
rect 17677 15058 17743 15061
rect 18469 15058 19269 15088
rect 17677 15056 19269 15058
rect 17677 15000 17682 15056
rect 17738 15000 19269 15056
rect 17677 14998 19269 15000
rect 12709 14995 12775 14996
rect 17677 14995 17743 14998
rect 18469 14968 19269 14998
rect 13813 14786 13879 14789
rect 14365 14788 14431 14789
rect 14365 14786 14412 14788
rect 13813 14784 14412 14786
rect 13813 14728 13818 14784
rect 13874 14728 14370 14784
rect 13813 14726 14412 14728
rect 13813 14723 13879 14726
rect 14365 14724 14412 14726
rect 14476 14724 14482 14788
rect 14365 14723 14431 14724
rect 3073 14720 3389 14721
rect 3073 14656 3079 14720
rect 3143 14656 3159 14720
rect 3223 14656 3239 14720
rect 3303 14656 3319 14720
rect 3383 14656 3389 14720
rect 3073 14655 3389 14656
rect 7328 14720 7644 14721
rect 7328 14656 7334 14720
rect 7398 14656 7414 14720
rect 7478 14656 7494 14720
rect 7558 14656 7574 14720
rect 7638 14656 7644 14720
rect 7328 14655 7644 14656
rect 11583 14720 11899 14721
rect 11583 14656 11589 14720
rect 11653 14656 11669 14720
rect 11733 14656 11749 14720
rect 11813 14656 11829 14720
rect 11893 14656 11899 14720
rect 11583 14655 11899 14656
rect 15838 14720 16154 14721
rect 15838 14656 15844 14720
rect 15908 14656 15924 14720
rect 15988 14656 16004 14720
rect 16068 14656 16084 14720
rect 16148 14656 16154 14720
rect 15838 14655 16154 14656
rect 841 14514 907 14517
rect 798 14512 907 14514
rect 798 14456 846 14512
rect 902 14456 907 14512
rect 798 14451 907 14456
rect 798 14408 858 14451
rect 0 14318 858 14408
rect 16941 14378 17007 14381
rect 18469 14378 19269 14408
rect 16941 14376 19269 14378
rect 16941 14320 16946 14376
rect 17002 14320 19269 14376
rect 16941 14318 19269 14320
rect 0 14288 800 14318
rect 16941 14315 17007 14318
rect 18469 14288 19269 14318
rect 3733 14176 4049 14177
rect 3733 14112 3739 14176
rect 3803 14112 3819 14176
rect 3883 14112 3899 14176
rect 3963 14112 3979 14176
rect 4043 14112 4049 14176
rect 3733 14111 4049 14112
rect 7988 14176 8304 14177
rect 7988 14112 7994 14176
rect 8058 14112 8074 14176
rect 8138 14112 8154 14176
rect 8218 14112 8234 14176
rect 8298 14112 8304 14176
rect 7988 14111 8304 14112
rect 12243 14176 12559 14177
rect 12243 14112 12249 14176
rect 12313 14112 12329 14176
rect 12393 14112 12409 14176
rect 12473 14112 12489 14176
rect 12553 14112 12559 14176
rect 12243 14111 12559 14112
rect 16498 14176 16814 14177
rect 16498 14112 16504 14176
rect 16568 14112 16584 14176
rect 16648 14112 16664 14176
rect 16728 14112 16744 14176
rect 16808 14112 16814 14176
rect 16498 14111 16814 14112
rect 8753 13834 8819 13837
rect 8710 13832 8819 13834
rect 8710 13776 8758 13832
rect 8814 13776 8819 13832
rect 8710 13771 8819 13776
rect 10726 13772 10732 13836
rect 10796 13834 10802 13836
rect 13721 13834 13787 13837
rect 10796 13832 13787 13834
rect 10796 13776 13726 13832
rect 13782 13776 13787 13832
rect 10796 13774 13787 13776
rect 10796 13772 10802 13774
rect 13721 13771 13787 13774
rect 3073 13632 3389 13633
rect 3073 13568 3079 13632
rect 3143 13568 3159 13632
rect 3223 13568 3239 13632
rect 3303 13568 3319 13632
rect 3383 13568 3389 13632
rect 3073 13567 3389 13568
rect 7328 13632 7644 13633
rect 7328 13568 7334 13632
rect 7398 13568 7414 13632
rect 7478 13568 7494 13632
rect 7558 13568 7574 13632
rect 7638 13568 7644 13632
rect 7328 13567 7644 13568
rect 5993 13426 6059 13429
rect 8710 13426 8770 13771
rect 11583 13632 11899 13633
rect 11583 13568 11589 13632
rect 11653 13568 11669 13632
rect 11733 13568 11749 13632
rect 11813 13568 11829 13632
rect 11893 13568 11899 13632
rect 11583 13567 11899 13568
rect 15838 13632 16154 13633
rect 15838 13568 15844 13632
rect 15908 13568 15924 13632
rect 15988 13568 16004 13632
rect 16068 13568 16084 13632
rect 16148 13568 16154 13632
rect 15838 13567 16154 13568
rect 10726 13426 10732 13428
rect 5993 13424 10732 13426
rect 5993 13368 5998 13424
rect 6054 13368 10732 13424
rect 5993 13366 10732 13368
rect 5993 13363 6059 13366
rect 10726 13364 10732 13366
rect 10796 13364 10802 13428
rect 3733 13088 4049 13089
rect 0 13018 800 13048
rect 3733 13024 3739 13088
rect 3803 13024 3819 13088
rect 3883 13024 3899 13088
rect 3963 13024 3979 13088
rect 4043 13024 4049 13088
rect 3733 13023 4049 13024
rect 7988 13088 8304 13089
rect 7988 13024 7994 13088
rect 8058 13024 8074 13088
rect 8138 13024 8154 13088
rect 8218 13024 8234 13088
rect 8298 13024 8304 13088
rect 7988 13023 8304 13024
rect 12243 13088 12559 13089
rect 12243 13024 12249 13088
rect 12313 13024 12329 13088
rect 12393 13024 12409 13088
rect 12473 13024 12489 13088
rect 12553 13024 12559 13088
rect 12243 13023 12559 13024
rect 16498 13088 16814 13089
rect 16498 13024 16504 13088
rect 16568 13024 16584 13088
rect 16648 13024 16664 13088
rect 16728 13024 16744 13088
rect 16808 13024 16814 13088
rect 16498 13023 16814 13024
rect 1025 13018 1091 13021
rect 0 13016 1091 13018
rect 0 12960 1030 13016
rect 1086 12960 1091 13016
rect 0 12958 1091 12960
rect 0 12928 800 12958
rect 1025 12955 1091 12958
rect 17677 13018 17743 13021
rect 18469 13018 19269 13048
rect 17677 13016 19269 13018
rect 17677 12960 17682 13016
rect 17738 12960 19269 13016
rect 17677 12958 19269 12960
rect 17677 12955 17743 12958
rect 18469 12928 19269 12958
rect 3073 12544 3389 12545
rect 3073 12480 3079 12544
rect 3143 12480 3159 12544
rect 3223 12480 3239 12544
rect 3303 12480 3319 12544
rect 3383 12480 3389 12544
rect 3073 12479 3389 12480
rect 7328 12544 7644 12545
rect 7328 12480 7334 12544
rect 7398 12480 7414 12544
rect 7478 12480 7494 12544
rect 7558 12480 7574 12544
rect 7638 12480 7644 12544
rect 7328 12479 7644 12480
rect 11583 12544 11899 12545
rect 11583 12480 11589 12544
rect 11653 12480 11669 12544
rect 11733 12480 11749 12544
rect 11813 12480 11829 12544
rect 11893 12480 11899 12544
rect 11583 12479 11899 12480
rect 15838 12544 16154 12545
rect 15838 12480 15844 12544
rect 15908 12480 15924 12544
rect 15988 12480 16004 12544
rect 16068 12480 16084 12544
rect 16148 12480 16154 12544
rect 15838 12479 16154 12480
rect 16297 12474 16363 12477
rect 16573 12474 16639 12477
rect 16297 12472 16639 12474
rect 16297 12416 16302 12472
rect 16358 12416 16578 12472
rect 16634 12416 16639 12472
rect 16297 12414 16639 12416
rect 16297 12411 16363 12414
rect 16573 12411 16639 12414
rect 0 12338 800 12368
rect 1301 12338 1367 12341
rect 0 12336 1367 12338
rect 0 12280 1306 12336
rect 1362 12280 1367 12336
rect 0 12278 1367 12280
rect 0 12248 800 12278
rect 1301 12275 1367 12278
rect 3733 12000 4049 12001
rect 3733 11936 3739 12000
rect 3803 11936 3819 12000
rect 3883 11936 3899 12000
rect 3963 11936 3979 12000
rect 4043 11936 4049 12000
rect 3733 11935 4049 11936
rect 7988 12000 8304 12001
rect 7988 11936 7994 12000
rect 8058 11936 8074 12000
rect 8138 11936 8154 12000
rect 8218 11936 8234 12000
rect 8298 11936 8304 12000
rect 7988 11935 8304 11936
rect 12243 12000 12559 12001
rect 12243 11936 12249 12000
rect 12313 11936 12329 12000
rect 12393 11936 12409 12000
rect 12473 11936 12489 12000
rect 12553 11936 12559 12000
rect 12243 11935 12559 11936
rect 16498 12000 16814 12001
rect 16498 11936 16504 12000
rect 16568 11936 16584 12000
rect 16648 11936 16664 12000
rect 16728 11936 16744 12000
rect 16808 11936 16814 12000
rect 16498 11935 16814 11936
rect 3073 11456 3389 11457
rect 3073 11392 3079 11456
rect 3143 11392 3159 11456
rect 3223 11392 3239 11456
rect 3303 11392 3319 11456
rect 3383 11392 3389 11456
rect 3073 11391 3389 11392
rect 7328 11456 7644 11457
rect 7328 11392 7334 11456
rect 7398 11392 7414 11456
rect 7478 11392 7494 11456
rect 7558 11392 7574 11456
rect 7638 11392 7644 11456
rect 7328 11391 7644 11392
rect 11583 11456 11899 11457
rect 11583 11392 11589 11456
rect 11653 11392 11669 11456
rect 11733 11392 11749 11456
rect 11813 11392 11829 11456
rect 11893 11392 11899 11456
rect 11583 11391 11899 11392
rect 15838 11456 16154 11457
rect 15838 11392 15844 11456
rect 15908 11392 15924 11456
rect 15988 11392 16004 11456
rect 16068 11392 16084 11456
rect 16148 11392 16154 11456
rect 15838 11391 16154 11392
rect 0 10978 800 11008
rect 1485 10978 1551 10981
rect 0 10976 1551 10978
rect 0 10920 1490 10976
rect 1546 10920 1551 10976
rect 0 10918 1551 10920
rect 0 10888 800 10918
rect 1485 10915 1551 10918
rect 3733 10912 4049 10913
rect 3733 10848 3739 10912
rect 3803 10848 3819 10912
rect 3883 10848 3899 10912
rect 3963 10848 3979 10912
rect 4043 10848 4049 10912
rect 3733 10847 4049 10848
rect 7988 10912 8304 10913
rect 7988 10848 7994 10912
rect 8058 10848 8074 10912
rect 8138 10848 8154 10912
rect 8218 10848 8234 10912
rect 8298 10848 8304 10912
rect 7988 10847 8304 10848
rect 12243 10912 12559 10913
rect 12243 10848 12249 10912
rect 12313 10848 12329 10912
rect 12393 10848 12409 10912
rect 12473 10848 12489 10912
rect 12553 10848 12559 10912
rect 12243 10847 12559 10848
rect 16498 10912 16814 10913
rect 16498 10848 16504 10912
rect 16568 10848 16584 10912
rect 16648 10848 16664 10912
rect 16728 10848 16744 10912
rect 16808 10848 16814 10912
rect 16498 10847 16814 10848
rect 10777 10844 10843 10845
rect 10726 10780 10732 10844
rect 10796 10842 10843 10844
rect 10796 10840 10888 10842
rect 10838 10784 10888 10840
rect 10796 10782 10888 10784
rect 10796 10780 10843 10782
rect 10777 10779 10843 10780
rect 3550 10644 3556 10708
rect 3620 10706 3626 10708
rect 9489 10706 9555 10709
rect 3620 10704 9555 10706
rect 3620 10648 9494 10704
rect 9550 10648 9555 10704
rect 3620 10646 9555 10648
rect 3620 10644 3626 10646
rect 9489 10643 9555 10646
rect 3073 10368 3389 10369
rect 0 10298 800 10328
rect 3073 10304 3079 10368
rect 3143 10304 3159 10368
rect 3223 10304 3239 10368
rect 3303 10304 3319 10368
rect 3383 10304 3389 10368
rect 3073 10303 3389 10304
rect 7328 10368 7644 10369
rect 7328 10304 7334 10368
rect 7398 10304 7414 10368
rect 7478 10304 7494 10368
rect 7558 10304 7574 10368
rect 7638 10304 7644 10368
rect 7328 10303 7644 10304
rect 11583 10368 11899 10369
rect 11583 10304 11589 10368
rect 11653 10304 11669 10368
rect 11733 10304 11749 10368
rect 11813 10304 11829 10368
rect 11893 10304 11899 10368
rect 11583 10303 11899 10304
rect 15838 10368 16154 10369
rect 15838 10304 15844 10368
rect 15908 10304 15924 10368
rect 15988 10304 16004 10368
rect 16068 10304 16084 10368
rect 16148 10304 16154 10368
rect 15838 10303 16154 10304
rect 1209 10298 1275 10301
rect 12801 10300 12867 10301
rect 0 10296 1275 10298
rect 0 10240 1214 10296
rect 1270 10240 1275 10296
rect 0 10238 1275 10240
rect 0 10208 800 10238
rect 1209 10235 1275 10238
rect 12750 10236 12756 10300
rect 12820 10298 12867 10300
rect 17677 10298 17743 10301
rect 18469 10298 19269 10328
rect 12820 10296 12912 10298
rect 12862 10240 12912 10296
rect 12820 10238 12912 10240
rect 17677 10296 19269 10298
rect 17677 10240 17682 10296
rect 17738 10240 19269 10296
rect 17677 10238 19269 10240
rect 12820 10236 12867 10238
rect 12801 10235 12867 10236
rect 17677 10235 17743 10238
rect 18469 10208 19269 10238
rect 13353 10026 13419 10029
rect 13905 10026 13971 10029
rect 15009 10026 15075 10029
rect 13353 10024 15075 10026
rect 13353 9968 13358 10024
rect 13414 9968 13910 10024
rect 13966 9968 15014 10024
rect 15070 9968 15075 10024
rect 13353 9966 15075 9968
rect 13353 9963 13419 9966
rect 13905 9963 13971 9966
rect 15009 9963 15075 9966
rect 3733 9824 4049 9825
rect 3733 9760 3739 9824
rect 3803 9760 3819 9824
rect 3883 9760 3899 9824
rect 3963 9760 3979 9824
rect 4043 9760 4049 9824
rect 3733 9759 4049 9760
rect 7988 9824 8304 9825
rect 7988 9760 7994 9824
rect 8058 9760 8074 9824
rect 8138 9760 8154 9824
rect 8218 9760 8234 9824
rect 8298 9760 8304 9824
rect 7988 9759 8304 9760
rect 12243 9824 12559 9825
rect 12243 9760 12249 9824
rect 12313 9760 12329 9824
rect 12393 9760 12409 9824
rect 12473 9760 12489 9824
rect 12553 9760 12559 9824
rect 12243 9759 12559 9760
rect 16498 9824 16814 9825
rect 16498 9760 16504 9824
rect 16568 9760 16584 9824
rect 16648 9760 16664 9824
rect 16728 9760 16744 9824
rect 16808 9760 16814 9824
rect 16498 9759 16814 9760
rect 0 9618 800 9648
rect 1853 9618 1919 9621
rect 0 9616 1919 9618
rect 0 9560 1858 9616
rect 1914 9560 1919 9616
rect 0 9558 1919 9560
rect 0 9528 800 9558
rect 1853 9555 1919 9558
rect 4521 9618 4587 9621
rect 10685 9618 10751 9621
rect 11697 9618 11763 9621
rect 4521 9616 11763 9618
rect 4521 9560 4526 9616
rect 4582 9560 10690 9616
rect 10746 9560 11702 9616
rect 11758 9560 11763 9616
rect 4521 9558 11763 9560
rect 4521 9555 4587 9558
rect 10685 9555 10751 9558
rect 11697 9555 11763 9558
rect 3073 9280 3389 9281
rect 3073 9216 3079 9280
rect 3143 9216 3159 9280
rect 3223 9216 3239 9280
rect 3303 9216 3319 9280
rect 3383 9216 3389 9280
rect 3073 9215 3389 9216
rect 7328 9280 7644 9281
rect 7328 9216 7334 9280
rect 7398 9216 7414 9280
rect 7478 9216 7494 9280
rect 7558 9216 7574 9280
rect 7638 9216 7644 9280
rect 7328 9215 7644 9216
rect 11583 9280 11899 9281
rect 11583 9216 11589 9280
rect 11653 9216 11669 9280
rect 11733 9216 11749 9280
rect 11813 9216 11829 9280
rect 11893 9216 11899 9280
rect 11583 9215 11899 9216
rect 15838 9280 16154 9281
rect 15838 9216 15844 9280
rect 15908 9216 15924 9280
rect 15988 9216 16004 9280
rect 16068 9216 16084 9280
rect 16148 9216 16154 9280
rect 15838 9215 16154 9216
rect 3733 8736 4049 8737
rect 3733 8672 3739 8736
rect 3803 8672 3819 8736
rect 3883 8672 3899 8736
rect 3963 8672 3979 8736
rect 4043 8672 4049 8736
rect 3733 8671 4049 8672
rect 7988 8736 8304 8737
rect 7988 8672 7994 8736
rect 8058 8672 8074 8736
rect 8138 8672 8154 8736
rect 8218 8672 8234 8736
rect 8298 8672 8304 8736
rect 7988 8671 8304 8672
rect 12243 8736 12559 8737
rect 12243 8672 12249 8736
rect 12313 8672 12329 8736
rect 12393 8672 12409 8736
rect 12473 8672 12489 8736
rect 12553 8672 12559 8736
rect 12243 8671 12559 8672
rect 16498 8736 16814 8737
rect 16498 8672 16504 8736
rect 16568 8672 16584 8736
rect 16648 8672 16664 8736
rect 16728 8672 16744 8736
rect 16808 8672 16814 8736
rect 16498 8671 16814 8672
rect 3601 8394 3667 8397
rect 11237 8394 11303 8397
rect 3601 8392 11303 8394
rect 3601 8336 3606 8392
rect 3662 8336 11242 8392
rect 11298 8336 11303 8392
rect 3601 8334 11303 8336
rect 3601 8331 3667 8334
rect 11237 8331 11303 8334
rect 16941 8258 17007 8261
rect 18469 8258 19269 8288
rect 16941 8256 19269 8258
rect 16941 8200 16946 8256
rect 17002 8200 19269 8256
rect 16941 8198 19269 8200
rect 16941 8195 17007 8198
rect 3073 8192 3389 8193
rect 3073 8128 3079 8192
rect 3143 8128 3159 8192
rect 3223 8128 3239 8192
rect 3303 8128 3319 8192
rect 3383 8128 3389 8192
rect 3073 8127 3389 8128
rect 7328 8192 7644 8193
rect 7328 8128 7334 8192
rect 7398 8128 7414 8192
rect 7478 8128 7494 8192
rect 7558 8128 7574 8192
rect 7638 8128 7644 8192
rect 7328 8127 7644 8128
rect 11583 8192 11899 8193
rect 11583 8128 11589 8192
rect 11653 8128 11669 8192
rect 11733 8128 11749 8192
rect 11813 8128 11829 8192
rect 11893 8128 11899 8192
rect 11583 8127 11899 8128
rect 15838 8192 16154 8193
rect 15838 8128 15844 8192
rect 15908 8128 15924 8192
rect 15988 8128 16004 8192
rect 16068 8128 16084 8192
rect 16148 8128 16154 8192
rect 18469 8168 19269 8198
rect 15838 8127 16154 8128
rect 7373 7986 7439 7989
rect 10726 7986 10732 7988
rect 7373 7984 10732 7986
rect 7373 7928 7378 7984
rect 7434 7928 10732 7984
rect 7373 7926 10732 7928
rect 7373 7923 7439 7926
rect 10726 7924 10732 7926
rect 10796 7986 10802 7988
rect 14365 7986 14431 7989
rect 10796 7984 14431 7986
rect 10796 7928 14370 7984
rect 14426 7928 14431 7984
rect 10796 7926 14431 7928
rect 10796 7924 10802 7926
rect 14365 7923 14431 7926
rect 12525 7850 12591 7853
rect 14549 7850 14615 7853
rect 12525 7848 14615 7850
rect 12525 7792 12530 7848
rect 12586 7792 14554 7848
rect 14610 7792 14615 7848
rect 12525 7790 14615 7792
rect 12525 7787 12591 7790
rect 14549 7787 14615 7790
rect 3733 7648 4049 7649
rect 3733 7584 3739 7648
rect 3803 7584 3819 7648
rect 3883 7584 3899 7648
rect 3963 7584 3979 7648
rect 4043 7584 4049 7648
rect 3733 7583 4049 7584
rect 7988 7648 8304 7649
rect 7988 7584 7994 7648
rect 8058 7584 8074 7648
rect 8138 7584 8154 7648
rect 8218 7584 8234 7648
rect 8298 7584 8304 7648
rect 7988 7583 8304 7584
rect 12243 7648 12559 7649
rect 12243 7584 12249 7648
rect 12313 7584 12329 7648
rect 12393 7584 12409 7648
rect 12473 7584 12489 7648
rect 12553 7584 12559 7648
rect 12243 7583 12559 7584
rect 16498 7648 16814 7649
rect 16498 7584 16504 7648
rect 16568 7584 16584 7648
rect 16648 7584 16664 7648
rect 16728 7584 16744 7648
rect 16808 7584 16814 7648
rect 16498 7583 16814 7584
rect 17769 7578 17835 7581
rect 18469 7578 19269 7608
rect 17769 7576 19269 7578
rect 17769 7520 17774 7576
rect 17830 7520 19269 7576
rect 17769 7518 19269 7520
rect 17769 7515 17835 7518
rect 18469 7488 19269 7518
rect 11973 7442 12039 7445
rect 14917 7442 14983 7445
rect 11973 7440 14983 7442
rect 11973 7384 11978 7440
rect 12034 7384 14922 7440
rect 14978 7384 14983 7440
rect 11973 7382 14983 7384
rect 11973 7379 12039 7382
rect 14917 7379 14983 7382
rect 3073 7104 3389 7105
rect 3073 7040 3079 7104
rect 3143 7040 3159 7104
rect 3223 7040 3239 7104
rect 3303 7040 3319 7104
rect 3383 7040 3389 7104
rect 3073 7039 3389 7040
rect 7328 7104 7644 7105
rect 7328 7040 7334 7104
rect 7398 7040 7414 7104
rect 7478 7040 7494 7104
rect 7558 7040 7574 7104
rect 7638 7040 7644 7104
rect 7328 7039 7644 7040
rect 11583 7104 11899 7105
rect 11583 7040 11589 7104
rect 11653 7040 11669 7104
rect 11733 7040 11749 7104
rect 11813 7040 11829 7104
rect 11893 7040 11899 7104
rect 11583 7039 11899 7040
rect 15838 7104 16154 7105
rect 15838 7040 15844 7104
rect 15908 7040 15924 7104
rect 15988 7040 16004 7104
rect 16068 7040 16084 7104
rect 16148 7040 16154 7104
rect 15838 7039 16154 7040
rect 4429 6898 4495 6901
rect 9489 6898 9555 6901
rect 4429 6896 9555 6898
rect 4429 6840 4434 6896
rect 4490 6840 9494 6896
rect 9550 6840 9555 6896
rect 4429 6838 9555 6840
rect 4429 6835 4495 6838
rect 9489 6835 9555 6838
rect 9949 6898 10015 6901
rect 14825 6898 14891 6901
rect 9949 6896 14891 6898
rect 9949 6840 9954 6896
rect 10010 6840 14830 6896
rect 14886 6840 14891 6896
rect 9949 6838 14891 6840
rect 9949 6835 10015 6838
rect 14825 6835 14891 6838
rect 17769 6898 17835 6901
rect 18469 6898 19269 6928
rect 17769 6896 19269 6898
rect 17769 6840 17774 6896
rect 17830 6840 19269 6896
rect 17769 6838 19269 6840
rect 17769 6835 17835 6838
rect 18469 6808 19269 6838
rect 4889 6762 4955 6765
rect 11881 6762 11947 6765
rect 4889 6760 11947 6762
rect 4889 6704 4894 6760
rect 4950 6704 11886 6760
rect 11942 6704 11947 6760
rect 4889 6702 11947 6704
rect 4889 6699 4955 6702
rect 11881 6699 11947 6702
rect 6085 6626 6151 6629
rect 7373 6626 7439 6629
rect 6085 6624 7439 6626
rect 6085 6568 6090 6624
rect 6146 6568 7378 6624
rect 7434 6568 7439 6624
rect 6085 6566 7439 6568
rect 6085 6563 6151 6566
rect 7373 6563 7439 6566
rect 3733 6560 4049 6561
rect 3733 6496 3739 6560
rect 3803 6496 3819 6560
rect 3883 6496 3899 6560
rect 3963 6496 3979 6560
rect 4043 6496 4049 6560
rect 3733 6495 4049 6496
rect 7988 6560 8304 6561
rect 7988 6496 7994 6560
rect 8058 6496 8074 6560
rect 8138 6496 8154 6560
rect 8218 6496 8234 6560
rect 8298 6496 8304 6560
rect 7988 6495 8304 6496
rect 12243 6560 12559 6561
rect 12243 6496 12249 6560
rect 12313 6496 12329 6560
rect 12393 6496 12409 6560
rect 12473 6496 12489 6560
rect 12553 6496 12559 6560
rect 12243 6495 12559 6496
rect 16498 6560 16814 6561
rect 16498 6496 16504 6560
rect 16568 6496 16584 6560
rect 16648 6496 16664 6560
rect 16728 6496 16744 6560
rect 16808 6496 16814 6560
rect 16498 6495 16814 6496
rect 11881 6354 11947 6357
rect 13997 6354 14063 6357
rect 11881 6352 14063 6354
rect 11881 6296 11886 6352
rect 11942 6296 14002 6352
rect 14058 6296 14063 6352
rect 11881 6294 14063 6296
rect 11881 6291 11947 6294
rect 13997 6291 14063 6294
rect 6177 6218 6243 6221
rect 7281 6218 7347 6221
rect 6177 6216 7347 6218
rect 6177 6160 6182 6216
rect 6238 6160 7286 6216
rect 7342 6160 7347 6216
rect 6177 6158 7347 6160
rect 6177 6155 6243 6158
rect 7281 6155 7347 6158
rect 17769 6218 17835 6221
rect 18469 6218 19269 6248
rect 17769 6216 19269 6218
rect 17769 6160 17774 6216
rect 17830 6160 19269 6216
rect 17769 6158 19269 6160
rect 17769 6155 17835 6158
rect 18469 6128 19269 6158
rect 3073 6016 3389 6017
rect 3073 5952 3079 6016
rect 3143 5952 3159 6016
rect 3223 5952 3239 6016
rect 3303 5952 3319 6016
rect 3383 5952 3389 6016
rect 3073 5951 3389 5952
rect 7328 6016 7644 6017
rect 7328 5952 7334 6016
rect 7398 5952 7414 6016
rect 7478 5952 7494 6016
rect 7558 5952 7574 6016
rect 7638 5952 7644 6016
rect 7328 5951 7644 5952
rect 11583 6016 11899 6017
rect 11583 5952 11589 6016
rect 11653 5952 11669 6016
rect 11733 5952 11749 6016
rect 11813 5952 11829 6016
rect 11893 5952 11899 6016
rect 11583 5951 11899 5952
rect 15838 6016 16154 6017
rect 15838 5952 15844 6016
rect 15908 5952 15924 6016
rect 15988 5952 16004 6016
rect 16068 5952 16084 6016
rect 16148 5952 16154 6016
rect 15838 5951 16154 5952
rect 14365 5812 14431 5813
rect 14365 5810 14412 5812
rect 14320 5808 14412 5810
rect 14320 5752 14370 5808
rect 14320 5750 14412 5752
rect 14365 5748 14412 5750
rect 14476 5748 14482 5812
rect 14365 5747 14431 5748
rect 6913 5674 6979 5677
rect 7189 5674 7255 5677
rect 11237 5674 11303 5677
rect 14457 5674 14523 5677
rect 6913 5672 14523 5674
rect 6913 5616 6918 5672
rect 6974 5616 7194 5672
rect 7250 5616 11242 5672
rect 11298 5616 14462 5672
rect 14518 5616 14523 5672
rect 6913 5614 14523 5616
rect 6913 5611 6979 5614
rect 7189 5611 7255 5614
rect 11237 5611 11303 5614
rect 14457 5611 14523 5614
rect 17677 5538 17743 5541
rect 18469 5538 19269 5568
rect 17677 5536 19269 5538
rect 17677 5480 17682 5536
rect 17738 5480 19269 5536
rect 17677 5478 19269 5480
rect 17677 5475 17743 5478
rect 3733 5472 4049 5473
rect 3733 5408 3739 5472
rect 3803 5408 3819 5472
rect 3883 5408 3899 5472
rect 3963 5408 3979 5472
rect 4043 5408 4049 5472
rect 3733 5407 4049 5408
rect 7988 5472 8304 5473
rect 7988 5408 7994 5472
rect 8058 5408 8074 5472
rect 8138 5408 8154 5472
rect 8218 5408 8234 5472
rect 8298 5408 8304 5472
rect 7988 5407 8304 5408
rect 12243 5472 12559 5473
rect 12243 5408 12249 5472
rect 12313 5408 12329 5472
rect 12393 5408 12409 5472
rect 12473 5408 12489 5472
rect 12553 5408 12559 5472
rect 12243 5407 12559 5408
rect 16498 5472 16814 5473
rect 16498 5408 16504 5472
rect 16568 5408 16584 5472
rect 16648 5408 16664 5472
rect 16728 5408 16744 5472
rect 16808 5408 16814 5472
rect 18469 5448 19269 5478
rect 16498 5407 16814 5408
rect 5349 5130 5415 5133
rect 7005 5130 7071 5133
rect 8017 5130 8083 5133
rect 5349 5128 8083 5130
rect 5349 5072 5354 5128
rect 5410 5072 7010 5128
rect 7066 5072 8022 5128
rect 8078 5072 8083 5128
rect 5349 5070 8083 5072
rect 5349 5067 5415 5070
rect 7005 5067 7071 5070
rect 8017 5067 8083 5070
rect 3073 4928 3389 4929
rect 3073 4864 3079 4928
rect 3143 4864 3159 4928
rect 3223 4864 3239 4928
rect 3303 4864 3319 4928
rect 3383 4864 3389 4928
rect 3073 4863 3389 4864
rect 7328 4928 7644 4929
rect 7328 4864 7334 4928
rect 7398 4864 7414 4928
rect 7478 4864 7494 4928
rect 7558 4864 7574 4928
rect 7638 4864 7644 4928
rect 7328 4863 7644 4864
rect 11583 4928 11899 4929
rect 11583 4864 11589 4928
rect 11653 4864 11669 4928
rect 11733 4864 11749 4928
rect 11813 4864 11829 4928
rect 11893 4864 11899 4928
rect 11583 4863 11899 4864
rect 15838 4928 16154 4929
rect 15838 4864 15844 4928
rect 15908 4864 15924 4928
rect 15988 4864 16004 4928
rect 16068 4864 16084 4928
rect 16148 4864 16154 4928
rect 15838 4863 16154 4864
rect 6545 4858 6611 4861
rect 6913 4858 6979 4861
rect 6545 4856 6979 4858
rect 6545 4800 6550 4856
rect 6606 4800 6918 4856
rect 6974 4800 6979 4856
rect 6545 4798 6979 4800
rect 6545 4795 6611 4798
rect 6913 4795 6979 4798
rect 17585 4858 17651 4861
rect 18469 4858 19269 4888
rect 17585 4856 19269 4858
rect 17585 4800 17590 4856
rect 17646 4800 19269 4856
rect 17585 4798 19269 4800
rect 17585 4795 17651 4798
rect 18469 4768 19269 4798
rect 5165 4722 5231 4725
rect 9029 4722 9095 4725
rect 5165 4720 9095 4722
rect 5165 4664 5170 4720
rect 5226 4664 9034 4720
rect 9090 4664 9095 4720
rect 5165 4662 9095 4664
rect 5165 4659 5231 4662
rect 9029 4659 9095 4662
rect 6821 4586 6887 4589
rect 7281 4586 7347 4589
rect 6821 4584 7347 4586
rect 6821 4528 6826 4584
rect 6882 4528 7286 4584
rect 7342 4528 7347 4584
rect 6821 4526 7347 4528
rect 6821 4523 6887 4526
rect 7281 4523 7347 4526
rect 3733 4384 4049 4385
rect 3733 4320 3739 4384
rect 3803 4320 3819 4384
rect 3883 4320 3899 4384
rect 3963 4320 3979 4384
rect 4043 4320 4049 4384
rect 3733 4319 4049 4320
rect 7988 4384 8304 4385
rect 7988 4320 7994 4384
rect 8058 4320 8074 4384
rect 8138 4320 8154 4384
rect 8218 4320 8234 4384
rect 8298 4320 8304 4384
rect 7988 4319 8304 4320
rect 12243 4384 12559 4385
rect 12243 4320 12249 4384
rect 12313 4320 12329 4384
rect 12393 4320 12409 4384
rect 12473 4320 12489 4384
rect 12553 4320 12559 4384
rect 12243 4319 12559 4320
rect 16498 4384 16814 4385
rect 16498 4320 16504 4384
rect 16568 4320 16584 4384
rect 16648 4320 16664 4384
rect 16728 4320 16744 4384
rect 16808 4320 16814 4384
rect 16498 4319 16814 4320
rect 3073 3840 3389 3841
rect 3073 3776 3079 3840
rect 3143 3776 3159 3840
rect 3223 3776 3239 3840
rect 3303 3776 3319 3840
rect 3383 3776 3389 3840
rect 3073 3775 3389 3776
rect 7328 3840 7644 3841
rect 7328 3776 7334 3840
rect 7398 3776 7414 3840
rect 7478 3776 7494 3840
rect 7558 3776 7574 3840
rect 7638 3776 7644 3840
rect 7328 3775 7644 3776
rect 11583 3840 11899 3841
rect 11583 3776 11589 3840
rect 11653 3776 11669 3840
rect 11733 3776 11749 3840
rect 11813 3776 11829 3840
rect 11893 3776 11899 3840
rect 11583 3775 11899 3776
rect 15838 3840 16154 3841
rect 15838 3776 15844 3840
rect 15908 3776 15924 3840
rect 15988 3776 16004 3840
rect 16068 3776 16084 3840
rect 16148 3776 16154 3840
rect 15838 3775 16154 3776
rect 17677 3498 17743 3501
rect 18469 3498 19269 3528
rect 17677 3496 19269 3498
rect 17677 3440 17682 3496
rect 17738 3440 19269 3496
rect 17677 3438 19269 3440
rect 17677 3435 17743 3438
rect 18469 3408 19269 3438
rect 3733 3296 4049 3297
rect 3733 3232 3739 3296
rect 3803 3232 3819 3296
rect 3883 3232 3899 3296
rect 3963 3232 3979 3296
rect 4043 3232 4049 3296
rect 3733 3231 4049 3232
rect 7988 3296 8304 3297
rect 7988 3232 7994 3296
rect 8058 3232 8074 3296
rect 8138 3232 8154 3296
rect 8218 3232 8234 3296
rect 8298 3232 8304 3296
rect 7988 3231 8304 3232
rect 12243 3296 12559 3297
rect 12243 3232 12249 3296
rect 12313 3232 12329 3296
rect 12393 3232 12409 3296
rect 12473 3232 12489 3296
rect 12553 3232 12559 3296
rect 12243 3231 12559 3232
rect 16498 3296 16814 3297
rect 16498 3232 16504 3296
rect 16568 3232 16584 3296
rect 16648 3232 16664 3296
rect 16728 3232 16744 3296
rect 16808 3232 16814 3296
rect 16498 3231 16814 3232
rect 10133 2954 10199 2957
rect 14641 2954 14707 2957
rect 10133 2952 14707 2954
rect 10133 2896 10138 2952
rect 10194 2896 14646 2952
rect 14702 2896 14707 2952
rect 10133 2894 14707 2896
rect 10133 2891 10199 2894
rect 14641 2891 14707 2894
rect 3073 2752 3389 2753
rect 3073 2688 3079 2752
rect 3143 2688 3159 2752
rect 3223 2688 3239 2752
rect 3303 2688 3319 2752
rect 3383 2688 3389 2752
rect 3073 2687 3389 2688
rect 7328 2752 7644 2753
rect 7328 2688 7334 2752
rect 7398 2688 7414 2752
rect 7478 2688 7494 2752
rect 7558 2688 7574 2752
rect 7638 2688 7644 2752
rect 7328 2687 7644 2688
rect 11583 2752 11899 2753
rect 11583 2688 11589 2752
rect 11653 2688 11669 2752
rect 11733 2688 11749 2752
rect 11813 2688 11829 2752
rect 11893 2688 11899 2752
rect 11583 2687 11899 2688
rect 15838 2752 16154 2753
rect 15838 2688 15844 2752
rect 15908 2688 15924 2752
rect 15988 2688 16004 2752
rect 16068 2688 16084 2752
rect 16148 2688 16154 2752
rect 15838 2687 16154 2688
rect 3733 2208 4049 2209
rect 3733 2144 3739 2208
rect 3803 2144 3819 2208
rect 3883 2144 3899 2208
rect 3963 2144 3979 2208
rect 4043 2144 4049 2208
rect 3733 2143 4049 2144
rect 7988 2208 8304 2209
rect 7988 2144 7994 2208
rect 8058 2144 8074 2208
rect 8138 2144 8154 2208
rect 8218 2144 8234 2208
rect 8298 2144 8304 2208
rect 7988 2143 8304 2144
rect 12243 2208 12559 2209
rect 12243 2144 12249 2208
rect 12313 2144 12329 2208
rect 12393 2144 12409 2208
rect 12473 2144 12489 2208
rect 12553 2144 12559 2208
rect 12243 2143 12559 2144
rect 16498 2208 16814 2209
rect 16498 2144 16504 2208
rect 16568 2144 16584 2208
rect 16648 2144 16664 2208
rect 16728 2144 16744 2208
rect 16808 2144 16814 2208
rect 16498 2143 16814 2144
<< via3 >>
rect 3079 19068 3143 19072
rect 3079 19012 3083 19068
rect 3083 19012 3139 19068
rect 3139 19012 3143 19068
rect 3079 19008 3143 19012
rect 3159 19068 3223 19072
rect 3159 19012 3163 19068
rect 3163 19012 3219 19068
rect 3219 19012 3223 19068
rect 3159 19008 3223 19012
rect 3239 19068 3303 19072
rect 3239 19012 3243 19068
rect 3243 19012 3299 19068
rect 3299 19012 3303 19068
rect 3239 19008 3303 19012
rect 3319 19068 3383 19072
rect 3319 19012 3323 19068
rect 3323 19012 3379 19068
rect 3379 19012 3383 19068
rect 3319 19008 3383 19012
rect 7334 19068 7398 19072
rect 7334 19012 7338 19068
rect 7338 19012 7394 19068
rect 7394 19012 7398 19068
rect 7334 19008 7398 19012
rect 7414 19068 7478 19072
rect 7414 19012 7418 19068
rect 7418 19012 7474 19068
rect 7474 19012 7478 19068
rect 7414 19008 7478 19012
rect 7494 19068 7558 19072
rect 7494 19012 7498 19068
rect 7498 19012 7554 19068
rect 7554 19012 7558 19068
rect 7494 19008 7558 19012
rect 7574 19068 7638 19072
rect 7574 19012 7578 19068
rect 7578 19012 7634 19068
rect 7634 19012 7638 19068
rect 7574 19008 7638 19012
rect 11589 19068 11653 19072
rect 11589 19012 11593 19068
rect 11593 19012 11649 19068
rect 11649 19012 11653 19068
rect 11589 19008 11653 19012
rect 11669 19068 11733 19072
rect 11669 19012 11673 19068
rect 11673 19012 11729 19068
rect 11729 19012 11733 19068
rect 11669 19008 11733 19012
rect 11749 19068 11813 19072
rect 11749 19012 11753 19068
rect 11753 19012 11809 19068
rect 11809 19012 11813 19068
rect 11749 19008 11813 19012
rect 11829 19068 11893 19072
rect 11829 19012 11833 19068
rect 11833 19012 11889 19068
rect 11889 19012 11893 19068
rect 11829 19008 11893 19012
rect 15844 19068 15908 19072
rect 15844 19012 15848 19068
rect 15848 19012 15904 19068
rect 15904 19012 15908 19068
rect 15844 19008 15908 19012
rect 15924 19068 15988 19072
rect 15924 19012 15928 19068
rect 15928 19012 15984 19068
rect 15984 19012 15988 19068
rect 15924 19008 15988 19012
rect 16004 19068 16068 19072
rect 16004 19012 16008 19068
rect 16008 19012 16064 19068
rect 16064 19012 16068 19068
rect 16004 19008 16068 19012
rect 16084 19068 16148 19072
rect 16084 19012 16088 19068
rect 16088 19012 16144 19068
rect 16144 19012 16148 19068
rect 16084 19008 16148 19012
rect 3739 18524 3803 18528
rect 3739 18468 3743 18524
rect 3743 18468 3799 18524
rect 3799 18468 3803 18524
rect 3739 18464 3803 18468
rect 3819 18524 3883 18528
rect 3819 18468 3823 18524
rect 3823 18468 3879 18524
rect 3879 18468 3883 18524
rect 3819 18464 3883 18468
rect 3899 18524 3963 18528
rect 3899 18468 3903 18524
rect 3903 18468 3959 18524
rect 3959 18468 3963 18524
rect 3899 18464 3963 18468
rect 3979 18524 4043 18528
rect 3979 18468 3983 18524
rect 3983 18468 4039 18524
rect 4039 18468 4043 18524
rect 3979 18464 4043 18468
rect 7994 18524 8058 18528
rect 7994 18468 7998 18524
rect 7998 18468 8054 18524
rect 8054 18468 8058 18524
rect 7994 18464 8058 18468
rect 8074 18524 8138 18528
rect 8074 18468 8078 18524
rect 8078 18468 8134 18524
rect 8134 18468 8138 18524
rect 8074 18464 8138 18468
rect 8154 18524 8218 18528
rect 8154 18468 8158 18524
rect 8158 18468 8214 18524
rect 8214 18468 8218 18524
rect 8154 18464 8218 18468
rect 8234 18524 8298 18528
rect 8234 18468 8238 18524
rect 8238 18468 8294 18524
rect 8294 18468 8298 18524
rect 8234 18464 8298 18468
rect 12249 18524 12313 18528
rect 12249 18468 12253 18524
rect 12253 18468 12309 18524
rect 12309 18468 12313 18524
rect 12249 18464 12313 18468
rect 12329 18524 12393 18528
rect 12329 18468 12333 18524
rect 12333 18468 12389 18524
rect 12389 18468 12393 18524
rect 12329 18464 12393 18468
rect 12409 18524 12473 18528
rect 12409 18468 12413 18524
rect 12413 18468 12469 18524
rect 12469 18468 12473 18524
rect 12409 18464 12473 18468
rect 12489 18524 12553 18528
rect 12489 18468 12493 18524
rect 12493 18468 12549 18524
rect 12549 18468 12553 18524
rect 12489 18464 12553 18468
rect 16504 18524 16568 18528
rect 16504 18468 16508 18524
rect 16508 18468 16564 18524
rect 16564 18468 16568 18524
rect 16504 18464 16568 18468
rect 16584 18524 16648 18528
rect 16584 18468 16588 18524
rect 16588 18468 16644 18524
rect 16644 18468 16648 18524
rect 16584 18464 16648 18468
rect 16664 18524 16728 18528
rect 16664 18468 16668 18524
rect 16668 18468 16724 18524
rect 16724 18468 16728 18524
rect 16664 18464 16728 18468
rect 16744 18524 16808 18528
rect 16744 18468 16748 18524
rect 16748 18468 16804 18524
rect 16804 18468 16808 18524
rect 16744 18464 16808 18468
rect 3079 17980 3143 17984
rect 3079 17924 3083 17980
rect 3083 17924 3139 17980
rect 3139 17924 3143 17980
rect 3079 17920 3143 17924
rect 3159 17980 3223 17984
rect 3159 17924 3163 17980
rect 3163 17924 3219 17980
rect 3219 17924 3223 17980
rect 3159 17920 3223 17924
rect 3239 17980 3303 17984
rect 3239 17924 3243 17980
rect 3243 17924 3299 17980
rect 3299 17924 3303 17980
rect 3239 17920 3303 17924
rect 3319 17980 3383 17984
rect 3319 17924 3323 17980
rect 3323 17924 3379 17980
rect 3379 17924 3383 17980
rect 3319 17920 3383 17924
rect 7334 17980 7398 17984
rect 7334 17924 7338 17980
rect 7338 17924 7394 17980
rect 7394 17924 7398 17980
rect 7334 17920 7398 17924
rect 7414 17980 7478 17984
rect 7414 17924 7418 17980
rect 7418 17924 7474 17980
rect 7474 17924 7478 17980
rect 7414 17920 7478 17924
rect 7494 17980 7558 17984
rect 7494 17924 7498 17980
rect 7498 17924 7554 17980
rect 7554 17924 7558 17980
rect 7494 17920 7558 17924
rect 7574 17980 7638 17984
rect 7574 17924 7578 17980
rect 7578 17924 7634 17980
rect 7634 17924 7638 17980
rect 7574 17920 7638 17924
rect 11589 17980 11653 17984
rect 11589 17924 11593 17980
rect 11593 17924 11649 17980
rect 11649 17924 11653 17980
rect 11589 17920 11653 17924
rect 11669 17980 11733 17984
rect 11669 17924 11673 17980
rect 11673 17924 11729 17980
rect 11729 17924 11733 17980
rect 11669 17920 11733 17924
rect 11749 17980 11813 17984
rect 11749 17924 11753 17980
rect 11753 17924 11809 17980
rect 11809 17924 11813 17980
rect 11749 17920 11813 17924
rect 11829 17980 11893 17984
rect 11829 17924 11833 17980
rect 11833 17924 11889 17980
rect 11889 17924 11893 17980
rect 11829 17920 11893 17924
rect 15844 17980 15908 17984
rect 15844 17924 15848 17980
rect 15848 17924 15904 17980
rect 15904 17924 15908 17980
rect 15844 17920 15908 17924
rect 15924 17980 15988 17984
rect 15924 17924 15928 17980
rect 15928 17924 15984 17980
rect 15984 17924 15988 17980
rect 15924 17920 15988 17924
rect 16004 17980 16068 17984
rect 16004 17924 16008 17980
rect 16008 17924 16064 17980
rect 16064 17924 16068 17980
rect 16004 17920 16068 17924
rect 16084 17980 16148 17984
rect 16084 17924 16088 17980
rect 16088 17924 16144 17980
rect 16144 17924 16148 17980
rect 16084 17920 16148 17924
rect 3556 17716 3620 17780
rect 3739 17436 3803 17440
rect 3739 17380 3743 17436
rect 3743 17380 3799 17436
rect 3799 17380 3803 17436
rect 3739 17376 3803 17380
rect 3819 17436 3883 17440
rect 3819 17380 3823 17436
rect 3823 17380 3879 17436
rect 3879 17380 3883 17436
rect 3819 17376 3883 17380
rect 3899 17436 3963 17440
rect 3899 17380 3903 17436
rect 3903 17380 3959 17436
rect 3959 17380 3963 17436
rect 3899 17376 3963 17380
rect 3979 17436 4043 17440
rect 3979 17380 3983 17436
rect 3983 17380 4039 17436
rect 4039 17380 4043 17436
rect 3979 17376 4043 17380
rect 7994 17436 8058 17440
rect 7994 17380 7998 17436
rect 7998 17380 8054 17436
rect 8054 17380 8058 17436
rect 7994 17376 8058 17380
rect 8074 17436 8138 17440
rect 8074 17380 8078 17436
rect 8078 17380 8134 17436
rect 8134 17380 8138 17436
rect 8074 17376 8138 17380
rect 8154 17436 8218 17440
rect 8154 17380 8158 17436
rect 8158 17380 8214 17436
rect 8214 17380 8218 17436
rect 8154 17376 8218 17380
rect 8234 17436 8298 17440
rect 8234 17380 8238 17436
rect 8238 17380 8294 17436
rect 8294 17380 8298 17436
rect 8234 17376 8298 17380
rect 12249 17436 12313 17440
rect 12249 17380 12253 17436
rect 12253 17380 12309 17436
rect 12309 17380 12313 17436
rect 12249 17376 12313 17380
rect 12329 17436 12393 17440
rect 12329 17380 12333 17436
rect 12333 17380 12389 17436
rect 12389 17380 12393 17436
rect 12329 17376 12393 17380
rect 12409 17436 12473 17440
rect 12409 17380 12413 17436
rect 12413 17380 12469 17436
rect 12469 17380 12473 17436
rect 12409 17376 12473 17380
rect 12489 17436 12553 17440
rect 12489 17380 12493 17436
rect 12493 17380 12549 17436
rect 12549 17380 12553 17436
rect 12489 17376 12553 17380
rect 16504 17436 16568 17440
rect 16504 17380 16508 17436
rect 16508 17380 16564 17436
rect 16564 17380 16568 17436
rect 16504 17376 16568 17380
rect 16584 17436 16648 17440
rect 16584 17380 16588 17436
rect 16588 17380 16644 17436
rect 16644 17380 16648 17436
rect 16584 17376 16648 17380
rect 16664 17436 16728 17440
rect 16664 17380 16668 17436
rect 16668 17380 16724 17436
rect 16724 17380 16728 17436
rect 16664 17376 16728 17380
rect 16744 17436 16808 17440
rect 16744 17380 16748 17436
rect 16748 17380 16804 17436
rect 16804 17380 16808 17436
rect 16744 17376 16808 17380
rect 3079 16892 3143 16896
rect 3079 16836 3083 16892
rect 3083 16836 3139 16892
rect 3139 16836 3143 16892
rect 3079 16832 3143 16836
rect 3159 16892 3223 16896
rect 3159 16836 3163 16892
rect 3163 16836 3219 16892
rect 3219 16836 3223 16892
rect 3159 16832 3223 16836
rect 3239 16892 3303 16896
rect 3239 16836 3243 16892
rect 3243 16836 3299 16892
rect 3299 16836 3303 16892
rect 3239 16832 3303 16836
rect 3319 16892 3383 16896
rect 3319 16836 3323 16892
rect 3323 16836 3379 16892
rect 3379 16836 3383 16892
rect 3319 16832 3383 16836
rect 7334 16892 7398 16896
rect 7334 16836 7338 16892
rect 7338 16836 7394 16892
rect 7394 16836 7398 16892
rect 7334 16832 7398 16836
rect 7414 16892 7478 16896
rect 7414 16836 7418 16892
rect 7418 16836 7474 16892
rect 7474 16836 7478 16892
rect 7414 16832 7478 16836
rect 7494 16892 7558 16896
rect 7494 16836 7498 16892
rect 7498 16836 7554 16892
rect 7554 16836 7558 16892
rect 7494 16832 7558 16836
rect 7574 16892 7638 16896
rect 7574 16836 7578 16892
rect 7578 16836 7634 16892
rect 7634 16836 7638 16892
rect 7574 16832 7638 16836
rect 11589 16892 11653 16896
rect 11589 16836 11593 16892
rect 11593 16836 11649 16892
rect 11649 16836 11653 16892
rect 11589 16832 11653 16836
rect 11669 16892 11733 16896
rect 11669 16836 11673 16892
rect 11673 16836 11729 16892
rect 11729 16836 11733 16892
rect 11669 16832 11733 16836
rect 11749 16892 11813 16896
rect 11749 16836 11753 16892
rect 11753 16836 11809 16892
rect 11809 16836 11813 16892
rect 11749 16832 11813 16836
rect 11829 16892 11893 16896
rect 11829 16836 11833 16892
rect 11833 16836 11889 16892
rect 11889 16836 11893 16892
rect 11829 16832 11893 16836
rect 15844 16892 15908 16896
rect 15844 16836 15848 16892
rect 15848 16836 15904 16892
rect 15904 16836 15908 16892
rect 15844 16832 15908 16836
rect 15924 16892 15988 16896
rect 15924 16836 15928 16892
rect 15928 16836 15984 16892
rect 15984 16836 15988 16892
rect 15924 16832 15988 16836
rect 16004 16892 16068 16896
rect 16004 16836 16008 16892
rect 16008 16836 16064 16892
rect 16064 16836 16068 16892
rect 16004 16832 16068 16836
rect 16084 16892 16148 16896
rect 16084 16836 16088 16892
rect 16088 16836 16144 16892
rect 16144 16836 16148 16892
rect 16084 16832 16148 16836
rect 3739 16348 3803 16352
rect 3739 16292 3743 16348
rect 3743 16292 3799 16348
rect 3799 16292 3803 16348
rect 3739 16288 3803 16292
rect 3819 16348 3883 16352
rect 3819 16292 3823 16348
rect 3823 16292 3879 16348
rect 3879 16292 3883 16348
rect 3819 16288 3883 16292
rect 3899 16348 3963 16352
rect 3899 16292 3903 16348
rect 3903 16292 3959 16348
rect 3959 16292 3963 16348
rect 3899 16288 3963 16292
rect 3979 16348 4043 16352
rect 3979 16292 3983 16348
rect 3983 16292 4039 16348
rect 4039 16292 4043 16348
rect 3979 16288 4043 16292
rect 7994 16348 8058 16352
rect 7994 16292 7998 16348
rect 7998 16292 8054 16348
rect 8054 16292 8058 16348
rect 7994 16288 8058 16292
rect 8074 16348 8138 16352
rect 8074 16292 8078 16348
rect 8078 16292 8134 16348
rect 8134 16292 8138 16348
rect 8074 16288 8138 16292
rect 8154 16348 8218 16352
rect 8154 16292 8158 16348
rect 8158 16292 8214 16348
rect 8214 16292 8218 16348
rect 8154 16288 8218 16292
rect 8234 16348 8298 16352
rect 8234 16292 8238 16348
rect 8238 16292 8294 16348
rect 8294 16292 8298 16348
rect 8234 16288 8298 16292
rect 12249 16348 12313 16352
rect 12249 16292 12253 16348
rect 12253 16292 12309 16348
rect 12309 16292 12313 16348
rect 12249 16288 12313 16292
rect 12329 16348 12393 16352
rect 12329 16292 12333 16348
rect 12333 16292 12389 16348
rect 12389 16292 12393 16348
rect 12329 16288 12393 16292
rect 12409 16348 12473 16352
rect 12409 16292 12413 16348
rect 12413 16292 12469 16348
rect 12469 16292 12473 16348
rect 12409 16288 12473 16292
rect 12489 16348 12553 16352
rect 12489 16292 12493 16348
rect 12493 16292 12549 16348
rect 12549 16292 12553 16348
rect 12489 16288 12553 16292
rect 16504 16348 16568 16352
rect 16504 16292 16508 16348
rect 16508 16292 16564 16348
rect 16564 16292 16568 16348
rect 16504 16288 16568 16292
rect 16584 16348 16648 16352
rect 16584 16292 16588 16348
rect 16588 16292 16644 16348
rect 16644 16292 16648 16348
rect 16584 16288 16648 16292
rect 16664 16348 16728 16352
rect 16664 16292 16668 16348
rect 16668 16292 16724 16348
rect 16724 16292 16728 16348
rect 16664 16288 16728 16292
rect 16744 16348 16808 16352
rect 16744 16292 16748 16348
rect 16748 16292 16804 16348
rect 16804 16292 16808 16348
rect 16744 16288 16808 16292
rect 3079 15804 3143 15808
rect 3079 15748 3083 15804
rect 3083 15748 3139 15804
rect 3139 15748 3143 15804
rect 3079 15744 3143 15748
rect 3159 15804 3223 15808
rect 3159 15748 3163 15804
rect 3163 15748 3219 15804
rect 3219 15748 3223 15804
rect 3159 15744 3223 15748
rect 3239 15804 3303 15808
rect 3239 15748 3243 15804
rect 3243 15748 3299 15804
rect 3299 15748 3303 15804
rect 3239 15744 3303 15748
rect 3319 15804 3383 15808
rect 3319 15748 3323 15804
rect 3323 15748 3379 15804
rect 3379 15748 3383 15804
rect 3319 15744 3383 15748
rect 7334 15804 7398 15808
rect 7334 15748 7338 15804
rect 7338 15748 7394 15804
rect 7394 15748 7398 15804
rect 7334 15744 7398 15748
rect 7414 15804 7478 15808
rect 7414 15748 7418 15804
rect 7418 15748 7474 15804
rect 7474 15748 7478 15804
rect 7414 15744 7478 15748
rect 7494 15804 7558 15808
rect 7494 15748 7498 15804
rect 7498 15748 7554 15804
rect 7554 15748 7558 15804
rect 7494 15744 7558 15748
rect 7574 15804 7638 15808
rect 7574 15748 7578 15804
rect 7578 15748 7634 15804
rect 7634 15748 7638 15804
rect 7574 15744 7638 15748
rect 11589 15804 11653 15808
rect 11589 15748 11593 15804
rect 11593 15748 11649 15804
rect 11649 15748 11653 15804
rect 11589 15744 11653 15748
rect 11669 15804 11733 15808
rect 11669 15748 11673 15804
rect 11673 15748 11729 15804
rect 11729 15748 11733 15804
rect 11669 15744 11733 15748
rect 11749 15804 11813 15808
rect 11749 15748 11753 15804
rect 11753 15748 11809 15804
rect 11809 15748 11813 15804
rect 11749 15744 11813 15748
rect 11829 15804 11893 15808
rect 11829 15748 11833 15804
rect 11833 15748 11889 15804
rect 11889 15748 11893 15804
rect 11829 15744 11893 15748
rect 15844 15804 15908 15808
rect 15844 15748 15848 15804
rect 15848 15748 15904 15804
rect 15904 15748 15908 15804
rect 15844 15744 15908 15748
rect 15924 15804 15988 15808
rect 15924 15748 15928 15804
rect 15928 15748 15984 15804
rect 15984 15748 15988 15804
rect 15924 15744 15988 15748
rect 16004 15804 16068 15808
rect 16004 15748 16008 15804
rect 16008 15748 16064 15804
rect 16064 15748 16068 15804
rect 16004 15744 16068 15748
rect 16084 15804 16148 15808
rect 16084 15748 16088 15804
rect 16088 15748 16144 15804
rect 16144 15748 16148 15804
rect 16084 15744 16148 15748
rect 3739 15260 3803 15264
rect 3739 15204 3743 15260
rect 3743 15204 3799 15260
rect 3799 15204 3803 15260
rect 3739 15200 3803 15204
rect 3819 15260 3883 15264
rect 3819 15204 3823 15260
rect 3823 15204 3879 15260
rect 3879 15204 3883 15260
rect 3819 15200 3883 15204
rect 3899 15260 3963 15264
rect 3899 15204 3903 15260
rect 3903 15204 3959 15260
rect 3959 15204 3963 15260
rect 3899 15200 3963 15204
rect 3979 15260 4043 15264
rect 3979 15204 3983 15260
rect 3983 15204 4039 15260
rect 4039 15204 4043 15260
rect 3979 15200 4043 15204
rect 7994 15260 8058 15264
rect 7994 15204 7998 15260
rect 7998 15204 8054 15260
rect 8054 15204 8058 15260
rect 7994 15200 8058 15204
rect 8074 15260 8138 15264
rect 8074 15204 8078 15260
rect 8078 15204 8134 15260
rect 8134 15204 8138 15260
rect 8074 15200 8138 15204
rect 8154 15260 8218 15264
rect 8154 15204 8158 15260
rect 8158 15204 8214 15260
rect 8214 15204 8218 15260
rect 8154 15200 8218 15204
rect 8234 15260 8298 15264
rect 8234 15204 8238 15260
rect 8238 15204 8294 15260
rect 8294 15204 8298 15260
rect 8234 15200 8298 15204
rect 12249 15260 12313 15264
rect 12249 15204 12253 15260
rect 12253 15204 12309 15260
rect 12309 15204 12313 15260
rect 12249 15200 12313 15204
rect 12329 15260 12393 15264
rect 12329 15204 12333 15260
rect 12333 15204 12389 15260
rect 12389 15204 12393 15260
rect 12329 15200 12393 15204
rect 12409 15260 12473 15264
rect 12409 15204 12413 15260
rect 12413 15204 12469 15260
rect 12469 15204 12473 15260
rect 12409 15200 12473 15204
rect 12489 15260 12553 15264
rect 12489 15204 12493 15260
rect 12493 15204 12549 15260
rect 12549 15204 12553 15260
rect 12489 15200 12553 15204
rect 16504 15260 16568 15264
rect 16504 15204 16508 15260
rect 16508 15204 16564 15260
rect 16564 15204 16568 15260
rect 16504 15200 16568 15204
rect 16584 15260 16648 15264
rect 16584 15204 16588 15260
rect 16588 15204 16644 15260
rect 16644 15204 16648 15260
rect 16584 15200 16648 15204
rect 16664 15260 16728 15264
rect 16664 15204 16668 15260
rect 16668 15204 16724 15260
rect 16724 15204 16728 15260
rect 16664 15200 16728 15204
rect 16744 15260 16808 15264
rect 16744 15204 16748 15260
rect 16748 15204 16804 15260
rect 16804 15204 16808 15260
rect 16744 15200 16808 15204
rect 12756 15056 12820 15060
rect 12756 15000 12770 15056
rect 12770 15000 12820 15056
rect 12756 14996 12820 15000
rect 14412 14784 14476 14788
rect 14412 14728 14426 14784
rect 14426 14728 14476 14784
rect 14412 14724 14476 14728
rect 3079 14716 3143 14720
rect 3079 14660 3083 14716
rect 3083 14660 3139 14716
rect 3139 14660 3143 14716
rect 3079 14656 3143 14660
rect 3159 14716 3223 14720
rect 3159 14660 3163 14716
rect 3163 14660 3219 14716
rect 3219 14660 3223 14716
rect 3159 14656 3223 14660
rect 3239 14716 3303 14720
rect 3239 14660 3243 14716
rect 3243 14660 3299 14716
rect 3299 14660 3303 14716
rect 3239 14656 3303 14660
rect 3319 14716 3383 14720
rect 3319 14660 3323 14716
rect 3323 14660 3379 14716
rect 3379 14660 3383 14716
rect 3319 14656 3383 14660
rect 7334 14716 7398 14720
rect 7334 14660 7338 14716
rect 7338 14660 7394 14716
rect 7394 14660 7398 14716
rect 7334 14656 7398 14660
rect 7414 14716 7478 14720
rect 7414 14660 7418 14716
rect 7418 14660 7474 14716
rect 7474 14660 7478 14716
rect 7414 14656 7478 14660
rect 7494 14716 7558 14720
rect 7494 14660 7498 14716
rect 7498 14660 7554 14716
rect 7554 14660 7558 14716
rect 7494 14656 7558 14660
rect 7574 14716 7638 14720
rect 7574 14660 7578 14716
rect 7578 14660 7634 14716
rect 7634 14660 7638 14716
rect 7574 14656 7638 14660
rect 11589 14716 11653 14720
rect 11589 14660 11593 14716
rect 11593 14660 11649 14716
rect 11649 14660 11653 14716
rect 11589 14656 11653 14660
rect 11669 14716 11733 14720
rect 11669 14660 11673 14716
rect 11673 14660 11729 14716
rect 11729 14660 11733 14716
rect 11669 14656 11733 14660
rect 11749 14716 11813 14720
rect 11749 14660 11753 14716
rect 11753 14660 11809 14716
rect 11809 14660 11813 14716
rect 11749 14656 11813 14660
rect 11829 14716 11893 14720
rect 11829 14660 11833 14716
rect 11833 14660 11889 14716
rect 11889 14660 11893 14716
rect 11829 14656 11893 14660
rect 15844 14716 15908 14720
rect 15844 14660 15848 14716
rect 15848 14660 15904 14716
rect 15904 14660 15908 14716
rect 15844 14656 15908 14660
rect 15924 14716 15988 14720
rect 15924 14660 15928 14716
rect 15928 14660 15984 14716
rect 15984 14660 15988 14716
rect 15924 14656 15988 14660
rect 16004 14716 16068 14720
rect 16004 14660 16008 14716
rect 16008 14660 16064 14716
rect 16064 14660 16068 14716
rect 16004 14656 16068 14660
rect 16084 14716 16148 14720
rect 16084 14660 16088 14716
rect 16088 14660 16144 14716
rect 16144 14660 16148 14716
rect 16084 14656 16148 14660
rect 3739 14172 3803 14176
rect 3739 14116 3743 14172
rect 3743 14116 3799 14172
rect 3799 14116 3803 14172
rect 3739 14112 3803 14116
rect 3819 14172 3883 14176
rect 3819 14116 3823 14172
rect 3823 14116 3879 14172
rect 3879 14116 3883 14172
rect 3819 14112 3883 14116
rect 3899 14172 3963 14176
rect 3899 14116 3903 14172
rect 3903 14116 3959 14172
rect 3959 14116 3963 14172
rect 3899 14112 3963 14116
rect 3979 14172 4043 14176
rect 3979 14116 3983 14172
rect 3983 14116 4039 14172
rect 4039 14116 4043 14172
rect 3979 14112 4043 14116
rect 7994 14172 8058 14176
rect 7994 14116 7998 14172
rect 7998 14116 8054 14172
rect 8054 14116 8058 14172
rect 7994 14112 8058 14116
rect 8074 14172 8138 14176
rect 8074 14116 8078 14172
rect 8078 14116 8134 14172
rect 8134 14116 8138 14172
rect 8074 14112 8138 14116
rect 8154 14172 8218 14176
rect 8154 14116 8158 14172
rect 8158 14116 8214 14172
rect 8214 14116 8218 14172
rect 8154 14112 8218 14116
rect 8234 14172 8298 14176
rect 8234 14116 8238 14172
rect 8238 14116 8294 14172
rect 8294 14116 8298 14172
rect 8234 14112 8298 14116
rect 12249 14172 12313 14176
rect 12249 14116 12253 14172
rect 12253 14116 12309 14172
rect 12309 14116 12313 14172
rect 12249 14112 12313 14116
rect 12329 14172 12393 14176
rect 12329 14116 12333 14172
rect 12333 14116 12389 14172
rect 12389 14116 12393 14172
rect 12329 14112 12393 14116
rect 12409 14172 12473 14176
rect 12409 14116 12413 14172
rect 12413 14116 12469 14172
rect 12469 14116 12473 14172
rect 12409 14112 12473 14116
rect 12489 14172 12553 14176
rect 12489 14116 12493 14172
rect 12493 14116 12549 14172
rect 12549 14116 12553 14172
rect 12489 14112 12553 14116
rect 16504 14172 16568 14176
rect 16504 14116 16508 14172
rect 16508 14116 16564 14172
rect 16564 14116 16568 14172
rect 16504 14112 16568 14116
rect 16584 14172 16648 14176
rect 16584 14116 16588 14172
rect 16588 14116 16644 14172
rect 16644 14116 16648 14172
rect 16584 14112 16648 14116
rect 16664 14172 16728 14176
rect 16664 14116 16668 14172
rect 16668 14116 16724 14172
rect 16724 14116 16728 14172
rect 16664 14112 16728 14116
rect 16744 14172 16808 14176
rect 16744 14116 16748 14172
rect 16748 14116 16804 14172
rect 16804 14116 16808 14172
rect 16744 14112 16808 14116
rect 10732 13772 10796 13836
rect 3079 13628 3143 13632
rect 3079 13572 3083 13628
rect 3083 13572 3139 13628
rect 3139 13572 3143 13628
rect 3079 13568 3143 13572
rect 3159 13628 3223 13632
rect 3159 13572 3163 13628
rect 3163 13572 3219 13628
rect 3219 13572 3223 13628
rect 3159 13568 3223 13572
rect 3239 13628 3303 13632
rect 3239 13572 3243 13628
rect 3243 13572 3299 13628
rect 3299 13572 3303 13628
rect 3239 13568 3303 13572
rect 3319 13628 3383 13632
rect 3319 13572 3323 13628
rect 3323 13572 3379 13628
rect 3379 13572 3383 13628
rect 3319 13568 3383 13572
rect 7334 13628 7398 13632
rect 7334 13572 7338 13628
rect 7338 13572 7394 13628
rect 7394 13572 7398 13628
rect 7334 13568 7398 13572
rect 7414 13628 7478 13632
rect 7414 13572 7418 13628
rect 7418 13572 7474 13628
rect 7474 13572 7478 13628
rect 7414 13568 7478 13572
rect 7494 13628 7558 13632
rect 7494 13572 7498 13628
rect 7498 13572 7554 13628
rect 7554 13572 7558 13628
rect 7494 13568 7558 13572
rect 7574 13628 7638 13632
rect 7574 13572 7578 13628
rect 7578 13572 7634 13628
rect 7634 13572 7638 13628
rect 7574 13568 7638 13572
rect 11589 13628 11653 13632
rect 11589 13572 11593 13628
rect 11593 13572 11649 13628
rect 11649 13572 11653 13628
rect 11589 13568 11653 13572
rect 11669 13628 11733 13632
rect 11669 13572 11673 13628
rect 11673 13572 11729 13628
rect 11729 13572 11733 13628
rect 11669 13568 11733 13572
rect 11749 13628 11813 13632
rect 11749 13572 11753 13628
rect 11753 13572 11809 13628
rect 11809 13572 11813 13628
rect 11749 13568 11813 13572
rect 11829 13628 11893 13632
rect 11829 13572 11833 13628
rect 11833 13572 11889 13628
rect 11889 13572 11893 13628
rect 11829 13568 11893 13572
rect 15844 13628 15908 13632
rect 15844 13572 15848 13628
rect 15848 13572 15904 13628
rect 15904 13572 15908 13628
rect 15844 13568 15908 13572
rect 15924 13628 15988 13632
rect 15924 13572 15928 13628
rect 15928 13572 15984 13628
rect 15984 13572 15988 13628
rect 15924 13568 15988 13572
rect 16004 13628 16068 13632
rect 16004 13572 16008 13628
rect 16008 13572 16064 13628
rect 16064 13572 16068 13628
rect 16004 13568 16068 13572
rect 16084 13628 16148 13632
rect 16084 13572 16088 13628
rect 16088 13572 16144 13628
rect 16144 13572 16148 13628
rect 16084 13568 16148 13572
rect 10732 13364 10796 13428
rect 3739 13084 3803 13088
rect 3739 13028 3743 13084
rect 3743 13028 3799 13084
rect 3799 13028 3803 13084
rect 3739 13024 3803 13028
rect 3819 13084 3883 13088
rect 3819 13028 3823 13084
rect 3823 13028 3879 13084
rect 3879 13028 3883 13084
rect 3819 13024 3883 13028
rect 3899 13084 3963 13088
rect 3899 13028 3903 13084
rect 3903 13028 3959 13084
rect 3959 13028 3963 13084
rect 3899 13024 3963 13028
rect 3979 13084 4043 13088
rect 3979 13028 3983 13084
rect 3983 13028 4039 13084
rect 4039 13028 4043 13084
rect 3979 13024 4043 13028
rect 7994 13084 8058 13088
rect 7994 13028 7998 13084
rect 7998 13028 8054 13084
rect 8054 13028 8058 13084
rect 7994 13024 8058 13028
rect 8074 13084 8138 13088
rect 8074 13028 8078 13084
rect 8078 13028 8134 13084
rect 8134 13028 8138 13084
rect 8074 13024 8138 13028
rect 8154 13084 8218 13088
rect 8154 13028 8158 13084
rect 8158 13028 8214 13084
rect 8214 13028 8218 13084
rect 8154 13024 8218 13028
rect 8234 13084 8298 13088
rect 8234 13028 8238 13084
rect 8238 13028 8294 13084
rect 8294 13028 8298 13084
rect 8234 13024 8298 13028
rect 12249 13084 12313 13088
rect 12249 13028 12253 13084
rect 12253 13028 12309 13084
rect 12309 13028 12313 13084
rect 12249 13024 12313 13028
rect 12329 13084 12393 13088
rect 12329 13028 12333 13084
rect 12333 13028 12389 13084
rect 12389 13028 12393 13084
rect 12329 13024 12393 13028
rect 12409 13084 12473 13088
rect 12409 13028 12413 13084
rect 12413 13028 12469 13084
rect 12469 13028 12473 13084
rect 12409 13024 12473 13028
rect 12489 13084 12553 13088
rect 12489 13028 12493 13084
rect 12493 13028 12549 13084
rect 12549 13028 12553 13084
rect 12489 13024 12553 13028
rect 16504 13084 16568 13088
rect 16504 13028 16508 13084
rect 16508 13028 16564 13084
rect 16564 13028 16568 13084
rect 16504 13024 16568 13028
rect 16584 13084 16648 13088
rect 16584 13028 16588 13084
rect 16588 13028 16644 13084
rect 16644 13028 16648 13084
rect 16584 13024 16648 13028
rect 16664 13084 16728 13088
rect 16664 13028 16668 13084
rect 16668 13028 16724 13084
rect 16724 13028 16728 13084
rect 16664 13024 16728 13028
rect 16744 13084 16808 13088
rect 16744 13028 16748 13084
rect 16748 13028 16804 13084
rect 16804 13028 16808 13084
rect 16744 13024 16808 13028
rect 3079 12540 3143 12544
rect 3079 12484 3083 12540
rect 3083 12484 3139 12540
rect 3139 12484 3143 12540
rect 3079 12480 3143 12484
rect 3159 12540 3223 12544
rect 3159 12484 3163 12540
rect 3163 12484 3219 12540
rect 3219 12484 3223 12540
rect 3159 12480 3223 12484
rect 3239 12540 3303 12544
rect 3239 12484 3243 12540
rect 3243 12484 3299 12540
rect 3299 12484 3303 12540
rect 3239 12480 3303 12484
rect 3319 12540 3383 12544
rect 3319 12484 3323 12540
rect 3323 12484 3379 12540
rect 3379 12484 3383 12540
rect 3319 12480 3383 12484
rect 7334 12540 7398 12544
rect 7334 12484 7338 12540
rect 7338 12484 7394 12540
rect 7394 12484 7398 12540
rect 7334 12480 7398 12484
rect 7414 12540 7478 12544
rect 7414 12484 7418 12540
rect 7418 12484 7474 12540
rect 7474 12484 7478 12540
rect 7414 12480 7478 12484
rect 7494 12540 7558 12544
rect 7494 12484 7498 12540
rect 7498 12484 7554 12540
rect 7554 12484 7558 12540
rect 7494 12480 7558 12484
rect 7574 12540 7638 12544
rect 7574 12484 7578 12540
rect 7578 12484 7634 12540
rect 7634 12484 7638 12540
rect 7574 12480 7638 12484
rect 11589 12540 11653 12544
rect 11589 12484 11593 12540
rect 11593 12484 11649 12540
rect 11649 12484 11653 12540
rect 11589 12480 11653 12484
rect 11669 12540 11733 12544
rect 11669 12484 11673 12540
rect 11673 12484 11729 12540
rect 11729 12484 11733 12540
rect 11669 12480 11733 12484
rect 11749 12540 11813 12544
rect 11749 12484 11753 12540
rect 11753 12484 11809 12540
rect 11809 12484 11813 12540
rect 11749 12480 11813 12484
rect 11829 12540 11893 12544
rect 11829 12484 11833 12540
rect 11833 12484 11889 12540
rect 11889 12484 11893 12540
rect 11829 12480 11893 12484
rect 15844 12540 15908 12544
rect 15844 12484 15848 12540
rect 15848 12484 15904 12540
rect 15904 12484 15908 12540
rect 15844 12480 15908 12484
rect 15924 12540 15988 12544
rect 15924 12484 15928 12540
rect 15928 12484 15984 12540
rect 15984 12484 15988 12540
rect 15924 12480 15988 12484
rect 16004 12540 16068 12544
rect 16004 12484 16008 12540
rect 16008 12484 16064 12540
rect 16064 12484 16068 12540
rect 16004 12480 16068 12484
rect 16084 12540 16148 12544
rect 16084 12484 16088 12540
rect 16088 12484 16144 12540
rect 16144 12484 16148 12540
rect 16084 12480 16148 12484
rect 3739 11996 3803 12000
rect 3739 11940 3743 11996
rect 3743 11940 3799 11996
rect 3799 11940 3803 11996
rect 3739 11936 3803 11940
rect 3819 11996 3883 12000
rect 3819 11940 3823 11996
rect 3823 11940 3879 11996
rect 3879 11940 3883 11996
rect 3819 11936 3883 11940
rect 3899 11996 3963 12000
rect 3899 11940 3903 11996
rect 3903 11940 3959 11996
rect 3959 11940 3963 11996
rect 3899 11936 3963 11940
rect 3979 11996 4043 12000
rect 3979 11940 3983 11996
rect 3983 11940 4039 11996
rect 4039 11940 4043 11996
rect 3979 11936 4043 11940
rect 7994 11996 8058 12000
rect 7994 11940 7998 11996
rect 7998 11940 8054 11996
rect 8054 11940 8058 11996
rect 7994 11936 8058 11940
rect 8074 11996 8138 12000
rect 8074 11940 8078 11996
rect 8078 11940 8134 11996
rect 8134 11940 8138 11996
rect 8074 11936 8138 11940
rect 8154 11996 8218 12000
rect 8154 11940 8158 11996
rect 8158 11940 8214 11996
rect 8214 11940 8218 11996
rect 8154 11936 8218 11940
rect 8234 11996 8298 12000
rect 8234 11940 8238 11996
rect 8238 11940 8294 11996
rect 8294 11940 8298 11996
rect 8234 11936 8298 11940
rect 12249 11996 12313 12000
rect 12249 11940 12253 11996
rect 12253 11940 12309 11996
rect 12309 11940 12313 11996
rect 12249 11936 12313 11940
rect 12329 11996 12393 12000
rect 12329 11940 12333 11996
rect 12333 11940 12389 11996
rect 12389 11940 12393 11996
rect 12329 11936 12393 11940
rect 12409 11996 12473 12000
rect 12409 11940 12413 11996
rect 12413 11940 12469 11996
rect 12469 11940 12473 11996
rect 12409 11936 12473 11940
rect 12489 11996 12553 12000
rect 12489 11940 12493 11996
rect 12493 11940 12549 11996
rect 12549 11940 12553 11996
rect 12489 11936 12553 11940
rect 16504 11996 16568 12000
rect 16504 11940 16508 11996
rect 16508 11940 16564 11996
rect 16564 11940 16568 11996
rect 16504 11936 16568 11940
rect 16584 11996 16648 12000
rect 16584 11940 16588 11996
rect 16588 11940 16644 11996
rect 16644 11940 16648 11996
rect 16584 11936 16648 11940
rect 16664 11996 16728 12000
rect 16664 11940 16668 11996
rect 16668 11940 16724 11996
rect 16724 11940 16728 11996
rect 16664 11936 16728 11940
rect 16744 11996 16808 12000
rect 16744 11940 16748 11996
rect 16748 11940 16804 11996
rect 16804 11940 16808 11996
rect 16744 11936 16808 11940
rect 3079 11452 3143 11456
rect 3079 11396 3083 11452
rect 3083 11396 3139 11452
rect 3139 11396 3143 11452
rect 3079 11392 3143 11396
rect 3159 11452 3223 11456
rect 3159 11396 3163 11452
rect 3163 11396 3219 11452
rect 3219 11396 3223 11452
rect 3159 11392 3223 11396
rect 3239 11452 3303 11456
rect 3239 11396 3243 11452
rect 3243 11396 3299 11452
rect 3299 11396 3303 11452
rect 3239 11392 3303 11396
rect 3319 11452 3383 11456
rect 3319 11396 3323 11452
rect 3323 11396 3379 11452
rect 3379 11396 3383 11452
rect 3319 11392 3383 11396
rect 7334 11452 7398 11456
rect 7334 11396 7338 11452
rect 7338 11396 7394 11452
rect 7394 11396 7398 11452
rect 7334 11392 7398 11396
rect 7414 11452 7478 11456
rect 7414 11396 7418 11452
rect 7418 11396 7474 11452
rect 7474 11396 7478 11452
rect 7414 11392 7478 11396
rect 7494 11452 7558 11456
rect 7494 11396 7498 11452
rect 7498 11396 7554 11452
rect 7554 11396 7558 11452
rect 7494 11392 7558 11396
rect 7574 11452 7638 11456
rect 7574 11396 7578 11452
rect 7578 11396 7634 11452
rect 7634 11396 7638 11452
rect 7574 11392 7638 11396
rect 11589 11452 11653 11456
rect 11589 11396 11593 11452
rect 11593 11396 11649 11452
rect 11649 11396 11653 11452
rect 11589 11392 11653 11396
rect 11669 11452 11733 11456
rect 11669 11396 11673 11452
rect 11673 11396 11729 11452
rect 11729 11396 11733 11452
rect 11669 11392 11733 11396
rect 11749 11452 11813 11456
rect 11749 11396 11753 11452
rect 11753 11396 11809 11452
rect 11809 11396 11813 11452
rect 11749 11392 11813 11396
rect 11829 11452 11893 11456
rect 11829 11396 11833 11452
rect 11833 11396 11889 11452
rect 11889 11396 11893 11452
rect 11829 11392 11893 11396
rect 15844 11452 15908 11456
rect 15844 11396 15848 11452
rect 15848 11396 15904 11452
rect 15904 11396 15908 11452
rect 15844 11392 15908 11396
rect 15924 11452 15988 11456
rect 15924 11396 15928 11452
rect 15928 11396 15984 11452
rect 15984 11396 15988 11452
rect 15924 11392 15988 11396
rect 16004 11452 16068 11456
rect 16004 11396 16008 11452
rect 16008 11396 16064 11452
rect 16064 11396 16068 11452
rect 16004 11392 16068 11396
rect 16084 11452 16148 11456
rect 16084 11396 16088 11452
rect 16088 11396 16144 11452
rect 16144 11396 16148 11452
rect 16084 11392 16148 11396
rect 3739 10908 3803 10912
rect 3739 10852 3743 10908
rect 3743 10852 3799 10908
rect 3799 10852 3803 10908
rect 3739 10848 3803 10852
rect 3819 10908 3883 10912
rect 3819 10852 3823 10908
rect 3823 10852 3879 10908
rect 3879 10852 3883 10908
rect 3819 10848 3883 10852
rect 3899 10908 3963 10912
rect 3899 10852 3903 10908
rect 3903 10852 3959 10908
rect 3959 10852 3963 10908
rect 3899 10848 3963 10852
rect 3979 10908 4043 10912
rect 3979 10852 3983 10908
rect 3983 10852 4039 10908
rect 4039 10852 4043 10908
rect 3979 10848 4043 10852
rect 7994 10908 8058 10912
rect 7994 10852 7998 10908
rect 7998 10852 8054 10908
rect 8054 10852 8058 10908
rect 7994 10848 8058 10852
rect 8074 10908 8138 10912
rect 8074 10852 8078 10908
rect 8078 10852 8134 10908
rect 8134 10852 8138 10908
rect 8074 10848 8138 10852
rect 8154 10908 8218 10912
rect 8154 10852 8158 10908
rect 8158 10852 8214 10908
rect 8214 10852 8218 10908
rect 8154 10848 8218 10852
rect 8234 10908 8298 10912
rect 8234 10852 8238 10908
rect 8238 10852 8294 10908
rect 8294 10852 8298 10908
rect 8234 10848 8298 10852
rect 12249 10908 12313 10912
rect 12249 10852 12253 10908
rect 12253 10852 12309 10908
rect 12309 10852 12313 10908
rect 12249 10848 12313 10852
rect 12329 10908 12393 10912
rect 12329 10852 12333 10908
rect 12333 10852 12389 10908
rect 12389 10852 12393 10908
rect 12329 10848 12393 10852
rect 12409 10908 12473 10912
rect 12409 10852 12413 10908
rect 12413 10852 12469 10908
rect 12469 10852 12473 10908
rect 12409 10848 12473 10852
rect 12489 10908 12553 10912
rect 12489 10852 12493 10908
rect 12493 10852 12549 10908
rect 12549 10852 12553 10908
rect 12489 10848 12553 10852
rect 16504 10908 16568 10912
rect 16504 10852 16508 10908
rect 16508 10852 16564 10908
rect 16564 10852 16568 10908
rect 16504 10848 16568 10852
rect 16584 10908 16648 10912
rect 16584 10852 16588 10908
rect 16588 10852 16644 10908
rect 16644 10852 16648 10908
rect 16584 10848 16648 10852
rect 16664 10908 16728 10912
rect 16664 10852 16668 10908
rect 16668 10852 16724 10908
rect 16724 10852 16728 10908
rect 16664 10848 16728 10852
rect 16744 10908 16808 10912
rect 16744 10852 16748 10908
rect 16748 10852 16804 10908
rect 16804 10852 16808 10908
rect 16744 10848 16808 10852
rect 10732 10840 10796 10844
rect 10732 10784 10782 10840
rect 10782 10784 10796 10840
rect 10732 10780 10796 10784
rect 3556 10644 3620 10708
rect 3079 10364 3143 10368
rect 3079 10308 3083 10364
rect 3083 10308 3139 10364
rect 3139 10308 3143 10364
rect 3079 10304 3143 10308
rect 3159 10364 3223 10368
rect 3159 10308 3163 10364
rect 3163 10308 3219 10364
rect 3219 10308 3223 10364
rect 3159 10304 3223 10308
rect 3239 10364 3303 10368
rect 3239 10308 3243 10364
rect 3243 10308 3299 10364
rect 3299 10308 3303 10364
rect 3239 10304 3303 10308
rect 3319 10364 3383 10368
rect 3319 10308 3323 10364
rect 3323 10308 3379 10364
rect 3379 10308 3383 10364
rect 3319 10304 3383 10308
rect 7334 10364 7398 10368
rect 7334 10308 7338 10364
rect 7338 10308 7394 10364
rect 7394 10308 7398 10364
rect 7334 10304 7398 10308
rect 7414 10364 7478 10368
rect 7414 10308 7418 10364
rect 7418 10308 7474 10364
rect 7474 10308 7478 10364
rect 7414 10304 7478 10308
rect 7494 10364 7558 10368
rect 7494 10308 7498 10364
rect 7498 10308 7554 10364
rect 7554 10308 7558 10364
rect 7494 10304 7558 10308
rect 7574 10364 7638 10368
rect 7574 10308 7578 10364
rect 7578 10308 7634 10364
rect 7634 10308 7638 10364
rect 7574 10304 7638 10308
rect 11589 10364 11653 10368
rect 11589 10308 11593 10364
rect 11593 10308 11649 10364
rect 11649 10308 11653 10364
rect 11589 10304 11653 10308
rect 11669 10364 11733 10368
rect 11669 10308 11673 10364
rect 11673 10308 11729 10364
rect 11729 10308 11733 10364
rect 11669 10304 11733 10308
rect 11749 10364 11813 10368
rect 11749 10308 11753 10364
rect 11753 10308 11809 10364
rect 11809 10308 11813 10364
rect 11749 10304 11813 10308
rect 11829 10364 11893 10368
rect 11829 10308 11833 10364
rect 11833 10308 11889 10364
rect 11889 10308 11893 10364
rect 11829 10304 11893 10308
rect 15844 10364 15908 10368
rect 15844 10308 15848 10364
rect 15848 10308 15904 10364
rect 15904 10308 15908 10364
rect 15844 10304 15908 10308
rect 15924 10364 15988 10368
rect 15924 10308 15928 10364
rect 15928 10308 15984 10364
rect 15984 10308 15988 10364
rect 15924 10304 15988 10308
rect 16004 10364 16068 10368
rect 16004 10308 16008 10364
rect 16008 10308 16064 10364
rect 16064 10308 16068 10364
rect 16004 10304 16068 10308
rect 16084 10364 16148 10368
rect 16084 10308 16088 10364
rect 16088 10308 16144 10364
rect 16144 10308 16148 10364
rect 16084 10304 16148 10308
rect 12756 10296 12820 10300
rect 12756 10240 12806 10296
rect 12806 10240 12820 10296
rect 12756 10236 12820 10240
rect 3739 9820 3803 9824
rect 3739 9764 3743 9820
rect 3743 9764 3799 9820
rect 3799 9764 3803 9820
rect 3739 9760 3803 9764
rect 3819 9820 3883 9824
rect 3819 9764 3823 9820
rect 3823 9764 3879 9820
rect 3879 9764 3883 9820
rect 3819 9760 3883 9764
rect 3899 9820 3963 9824
rect 3899 9764 3903 9820
rect 3903 9764 3959 9820
rect 3959 9764 3963 9820
rect 3899 9760 3963 9764
rect 3979 9820 4043 9824
rect 3979 9764 3983 9820
rect 3983 9764 4039 9820
rect 4039 9764 4043 9820
rect 3979 9760 4043 9764
rect 7994 9820 8058 9824
rect 7994 9764 7998 9820
rect 7998 9764 8054 9820
rect 8054 9764 8058 9820
rect 7994 9760 8058 9764
rect 8074 9820 8138 9824
rect 8074 9764 8078 9820
rect 8078 9764 8134 9820
rect 8134 9764 8138 9820
rect 8074 9760 8138 9764
rect 8154 9820 8218 9824
rect 8154 9764 8158 9820
rect 8158 9764 8214 9820
rect 8214 9764 8218 9820
rect 8154 9760 8218 9764
rect 8234 9820 8298 9824
rect 8234 9764 8238 9820
rect 8238 9764 8294 9820
rect 8294 9764 8298 9820
rect 8234 9760 8298 9764
rect 12249 9820 12313 9824
rect 12249 9764 12253 9820
rect 12253 9764 12309 9820
rect 12309 9764 12313 9820
rect 12249 9760 12313 9764
rect 12329 9820 12393 9824
rect 12329 9764 12333 9820
rect 12333 9764 12389 9820
rect 12389 9764 12393 9820
rect 12329 9760 12393 9764
rect 12409 9820 12473 9824
rect 12409 9764 12413 9820
rect 12413 9764 12469 9820
rect 12469 9764 12473 9820
rect 12409 9760 12473 9764
rect 12489 9820 12553 9824
rect 12489 9764 12493 9820
rect 12493 9764 12549 9820
rect 12549 9764 12553 9820
rect 12489 9760 12553 9764
rect 16504 9820 16568 9824
rect 16504 9764 16508 9820
rect 16508 9764 16564 9820
rect 16564 9764 16568 9820
rect 16504 9760 16568 9764
rect 16584 9820 16648 9824
rect 16584 9764 16588 9820
rect 16588 9764 16644 9820
rect 16644 9764 16648 9820
rect 16584 9760 16648 9764
rect 16664 9820 16728 9824
rect 16664 9764 16668 9820
rect 16668 9764 16724 9820
rect 16724 9764 16728 9820
rect 16664 9760 16728 9764
rect 16744 9820 16808 9824
rect 16744 9764 16748 9820
rect 16748 9764 16804 9820
rect 16804 9764 16808 9820
rect 16744 9760 16808 9764
rect 3079 9276 3143 9280
rect 3079 9220 3083 9276
rect 3083 9220 3139 9276
rect 3139 9220 3143 9276
rect 3079 9216 3143 9220
rect 3159 9276 3223 9280
rect 3159 9220 3163 9276
rect 3163 9220 3219 9276
rect 3219 9220 3223 9276
rect 3159 9216 3223 9220
rect 3239 9276 3303 9280
rect 3239 9220 3243 9276
rect 3243 9220 3299 9276
rect 3299 9220 3303 9276
rect 3239 9216 3303 9220
rect 3319 9276 3383 9280
rect 3319 9220 3323 9276
rect 3323 9220 3379 9276
rect 3379 9220 3383 9276
rect 3319 9216 3383 9220
rect 7334 9276 7398 9280
rect 7334 9220 7338 9276
rect 7338 9220 7394 9276
rect 7394 9220 7398 9276
rect 7334 9216 7398 9220
rect 7414 9276 7478 9280
rect 7414 9220 7418 9276
rect 7418 9220 7474 9276
rect 7474 9220 7478 9276
rect 7414 9216 7478 9220
rect 7494 9276 7558 9280
rect 7494 9220 7498 9276
rect 7498 9220 7554 9276
rect 7554 9220 7558 9276
rect 7494 9216 7558 9220
rect 7574 9276 7638 9280
rect 7574 9220 7578 9276
rect 7578 9220 7634 9276
rect 7634 9220 7638 9276
rect 7574 9216 7638 9220
rect 11589 9276 11653 9280
rect 11589 9220 11593 9276
rect 11593 9220 11649 9276
rect 11649 9220 11653 9276
rect 11589 9216 11653 9220
rect 11669 9276 11733 9280
rect 11669 9220 11673 9276
rect 11673 9220 11729 9276
rect 11729 9220 11733 9276
rect 11669 9216 11733 9220
rect 11749 9276 11813 9280
rect 11749 9220 11753 9276
rect 11753 9220 11809 9276
rect 11809 9220 11813 9276
rect 11749 9216 11813 9220
rect 11829 9276 11893 9280
rect 11829 9220 11833 9276
rect 11833 9220 11889 9276
rect 11889 9220 11893 9276
rect 11829 9216 11893 9220
rect 15844 9276 15908 9280
rect 15844 9220 15848 9276
rect 15848 9220 15904 9276
rect 15904 9220 15908 9276
rect 15844 9216 15908 9220
rect 15924 9276 15988 9280
rect 15924 9220 15928 9276
rect 15928 9220 15984 9276
rect 15984 9220 15988 9276
rect 15924 9216 15988 9220
rect 16004 9276 16068 9280
rect 16004 9220 16008 9276
rect 16008 9220 16064 9276
rect 16064 9220 16068 9276
rect 16004 9216 16068 9220
rect 16084 9276 16148 9280
rect 16084 9220 16088 9276
rect 16088 9220 16144 9276
rect 16144 9220 16148 9276
rect 16084 9216 16148 9220
rect 3739 8732 3803 8736
rect 3739 8676 3743 8732
rect 3743 8676 3799 8732
rect 3799 8676 3803 8732
rect 3739 8672 3803 8676
rect 3819 8732 3883 8736
rect 3819 8676 3823 8732
rect 3823 8676 3879 8732
rect 3879 8676 3883 8732
rect 3819 8672 3883 8676
rect 3899 8732 3963 8736
rect 3899 8676 3903 8732
rect 3903 8676 3959 8732
rect 3959 8676 3963 8732
rect 3899 8672 3963 8676
rect 3979 8732 4043 8736
rect 3979 8676 3983 8732
rect 3983 8676 4039 8732
rect 4039 8676 4043 8732
rect 3979 8672 4043 8676
rect 7994 8732 8058 8736
rect 7994 8676 7998 8732
rect 7998 8676 8054 8732
rect 8054 8676 8058 8732
rect 7994 8672 8058 8676
rect 8074 8732 8138 8736
rect 8074 8676 8078 8732
rect 8078 8676 8134 8732
rect 8134 8676 8138 8732
rect 8074 8672 8138 8676
rect 8154 8732 8218 8736
rect 8154 8676 8158 8732
rect 8158 8676 8214 8732
rect 8214 8676 8218 8732
rect 8154 8672 8218 8676
rect 8234 8732 8298 8736
rect 8234 8676 8238 8732
rect 8238 8676 8294 8732
rect 8294 8676 8298 8732
rect 8234 8672 8298 8676
rect 12249 8732 12313 8736
rect 12249 8676 12253 8732
rect 12253 8676 12309 8732
rect 12309 8676 12313 8732
rect 12249 8672 12313 8676
rect 12329 8732 12393 8736
rect 12329 8676 12333 8732
rect 12333 8676 12389 8732
rect 12389 8676 12393 8732
rect 12329 8672 12393 8676
rect 12409 8732 12473 8736
rect 12409 8676 12413 8732
rect 12413 8676 12469 8732
rect 12469 8676 12473 8732
rect 12409 8672 12473 8676
rect 12489 8732 12553 8736
rect 12489 8676 12493 8732
rect 12493 8676 12549 8732
rect 12549 8676 12553 8732
rect 12489 8672 12553 8676
rect 16504 8732 16568 8736
rect 16504 8676 16508 8732
rect 16508 8676 16564 8732
rect 16564 8676 16568 8732
rect 16504 8672 16568 8676
rect 16584 8732 16648 8736
rect 16584 8676 16588 8732
rect 16588 8676 16644 8732
rect 16644 8676 16648 8732
rect 16584 8672 16648 8676
rect 16664 8732 16728 8736
rect 16664 8676 16668 8732
rect 16668 8676 16724 8732
rect 16724 8676 16728 8732
rect 16664 8672 16728 8676
rect 16744 8732 16808 8736
rect 16744 8676 16748 8732
rect 16748 8676 16804 8732
rect 16804 8676 16808 8732
rect 16744 8672 16808 8676
rect 3079 8188 3143 8192
rect 3079 8132 3083 8188
rect 3083 8132 3139 8188
rect 3139 8132 3143 8188
rect 3079 8128 3143 8132
rect 3159 8188 3223 8192
rect 3159 8132 3163 8188
rect 3163 8132 3219 8188
rect 3219 8132 3223 8188
rect 3159 8128 3223 8132
rect 3239 8188 3303 8192
rect 3239 8132 3243 8188
rect 3243 8132 3299 8188
rect 3299 8132 3303 8188
rect 3239 8128 3303 8132
rect 3319 8188 3383 8192
rect 3319 8132 3323 8188
rect 3323 8132 3379 8188
rect 3379 8132 3383 8188
rect 3319 8128 3383 8132
rect 7334 8188 7398 8192
rect 7334 8132 7338 8188
rect 7338 8132 7394 8188
rect 7394 8132 7398 8188
rect 7334 8128 7398 8132
rect 7414 8188 7478 8192
rect 7414 8132 7418 8188
rect 7418 8132 7474 8188
rect 7474 8132 7478 8188
rect 7414 8128 7478 8132
rect 7494 8188 7558 8192
rect 7494 8132 7498 8188
rect 7498 8132 7554 8188
rect 7554 8132 7558 8188
rect 7494 8128 7558 8132
rect 7574 8188 7638 8192
rect 7574 8132 7578 8188
rect 7578 8132 7634 8188
rect 7634 8132 7638 8188
rect 7574 8128 7638 8132
rect 11589 8188 11653 8192
rect 11589 8132 11593 8188
rect 11593 8132 11649 8188
rect 11649 8132 11653 8188
rect 11589 8128 11653 8132
rect 11669 8188 11733 8192
rect 11669 8132 11673 8188
rect 11673 8132 11729 8188
rect 11729 8132 11733 8188
rect 11669 8128 11733 8132
rect 11749 8188 11813 8192
rect 11749 8132 11753 8188
rect 11753 8132 11809 8188
rect 11809 8132 11813 8188
rect 11749 8128 11813 8132
rect 11829 8188 11893 8192
rect 11829 8132 11833 8188
rect 11833 8132 11889 8188
rect 11889 8132 11893 8188
rect 11829 8128 11893 8132
rect 15844 8188 15908 8192
rect 15844 8132 15848 8188
rect 15848 8132 15904 8188
rect 15904 8132 15908 8188
rect 15844 8128 15908 8132
rect 15924 8188 15988 8192
rect 15924 8132 15928 8188
rect 15928 8132 15984 8188
rect 15984 8132 15988 8188
rect 15924 8128 15988 8132
rect 16004 8188 16068 8192
rect 16004 8132 16008 8188
rect 16008 8132 16064 8188
rect 16064 8132 16068 8188
rect 16004 8128 16068 8132
rect 16084 8188 16148 8192
rect 16084 8132 16088 8188
rect 16088 8132 16144 8188
rect 16144 8132 16148 8188
rect 16084 8128 16148 8132
rect 10732 7924 10796 7988
rect 3739 7644 3803 7648
rect 3739 7588 3743 7644
rect 3743 7588 3799 7644
rect 3799 7588 3803 7644
rect 3739 7584 3803 7588
rect 3819 7644 3883 7648
rect 3819 7588 3823 7644
rect 3823 7588 3879 7644
rect 3879 7588 3883 7644
rect 3819 7584 3883 7588
rect 3899 7644 3963 7648
rect 3899 7588 3903 7644
rect 3903 7588 3959 7644
rect 3959 7588 3963 7644
rect 3899 7584 3963 7588
rect 3979 7644 4043 7648
rect 3979 7588 3983 7644
rect 3983 7588 4039 7644
rect 4039 7588 4043 7644
rect 3979 7584 4043 7588
rect 7994 7644 8058 7648
rect 7994 7588 7998 7644
rect 7998 7588 8054 7644
rect 8054 7588 8058 7644
rect 7994 7584 8058 7588
rect 8074 7644 8138 7648
rect 8074 7588 8078 7644
rect 8078 7588 8134 7644
rect 8134 7588 8138 7644
rect 8074 7584 8138 7588
rect 8154 7644 8218 7648
rect 8154 7588 8158 7644
rect 8158 7588 8214 7644
rect 8214 7588 8218 7644
rect 8154 7584 8218 7588
rect 8234 7644 8298 7648
rect 8234 7588 8238 7644
rect 8238 7588 8294 7644
rect 8294 7588 8298 7644
rect 8234 7584 8298 7588
rect 12249 7644 12313 7648
rect 12249 7588 12253 7644
rect 12253 7588 12309 7644
rect 12309 7588 12313 7644
rect 12249 7584 12313 7588
rect 12329 7644 12393 7648
rect 12329 7588 12333 7644
rect 12333 7588 12389 7644
rect 12389 7588 12393 7644
rect 12329 7584 12393 7588
rect 12409 7644 12473 7648
rect 12409 7588 12413 7644
rect 12413 7588 12469 7644
rect 12469 7588 12473 7644
rect 12409 7584 12473 7588
rect 12489 7644 12553 7648
rect 12489 7588 12493 7644
rect 12493 7588 12549 7644
rect 12549 7588 12553 7644
rect 12489 7584 12553 7588
rect 16504 7644 16568 7648
rect 16504 7588 16508 7644
rect 16508 7588 16564 7644
rect 16564 7588 16568 7644
rect 16504 7584 16568 7588
rect 16584 7644 16648 7648
rect 16584 7588 16588 7644
rect 16588 7588 16644 7644
rect 16644 7588 16648 7644
rect 16584 7584 16648 7588
rect 16664 7644 16728 7648
rect 16664 7588 16668 7644
rect 16668 7588 16724 7644
rect 16724 7588 16728 7644
rect 16664 7584 16728 7588
rect 16744 7644 16808 7648
rect 16744 7588 16748 7644
rect 16748 7588 16804 7644
rect 16804 7588 16808 7644
rect 16744 7584 16808 7588
rect 3079 7100 3143 7104
rect 3079 7044 3083 7100
rect 3083 7044 3139 7100
rect 3139 7044 3143 7100
rect 3079 7040 3143 7044
rect 3159 7100 3223 7104
rect 3159 7044 3163 7100
rect 3163 7044 3219 7100
rect 3219 7044 3223 7100
rect 3159 7040 3223 7044
rect 3239 7100 3303 7104
rect 3239 7044 3243 7100
rect 3243 7044 3299 7100
rect 3299 7044 3303 7100
rect 3239 7040 3303 7044
rect 3319 7100 3383 7104
rect 3319 7044 3323 7100
rect 3323 7044 3379 7100
rect 3379 7044 3383 7100
rect 3319 7040 3383 7044
rect 7334 7100 7398 7104
rect 7334 7044 7338 7100
rect 7338 7044 7394 7100
rect 7394 7044 7398 7100
rect 7334 7040 7398 7044
rect 7414 7100 7478 7104
rect 7414 7044 7418 7100
rect 7418 7044 7474 7100
rect 7474 7044 7478 7100
rect 7414 7040 7478 7044
rect 7494 7100 7558 7104
rect 7494 7044 7498 7100
rect 7498 7044 7554 7100
rect 7554 7044 7558 7100
rect 7494 7040 7558 7044
rect 7574 7100 7638 7104
rect 7574 7044 7578 7100
rect 7578 7044 7634 7100
rect 7634 7044 7638 7100
rect 7574 7040 7638 7044
rect 11589 7100 11653 7104
rect 11589 7044 11593 7100
rect 11593 7044 11649 7100
rect 11649 7044 11653 7100
rect 11589 7040 11653 7044
rect 11669 7100 11733 7104
rect 11669 7044 11673 7100
rect 11673 7044 11729 7100
rect 11729 7044 11733 7100
rect 11669 7040 11733 7044
rect 11749 7100 11813 7104
rect 11749 7044 11753 7100
rect 11753 7044 11809 7100
rect 11809 7044 11813 7100
rect 11749 7040 11813 7044
rect 11829 7100 11893 7104
rect 11829 7044 11833 7100
rect 11833 7044 11889 7100
rect 11889 7044 11893 7100
rect 11829 7040 11893 7044
rect 15844 7100 15908 7104
rect 15844 7044 15848 7100
rect 15848 7044 15904 7100
rect 15904 7044 15908 7100
rect 15844 7040 15908 7044
rect 15924 7100 15988 7104
rect 15924 7044 15928 7100
rect 15928 7044 15984 7100
rect 15984 7044 15988 7100
rect 15924 7040 15988 7044
rect 16004 7100 16068 7104
rect 16004 7044 16008 7100
rect 16008 7044 16064 7100
rect 16064 7044 16068 7100
rect 16004 7040 16068 7044
rect 16084 7100 16148 7104
rect 16084 7044 16088 7100
rect 16088 7044 16144 7100
rect 16144 7044 16148 7100
rect 16084 7040 16148 7044
rect 3739 6556 3803 6560
rect 3739 6500 3743 6556
rect 3743 6500 3799 6556
rect 3799 6500 3803 6556
rect 3739 6496 3803 6500
rect 3819 6556 3883 6560
rect 3819 6500 3823 6556
rect 3823 6500 3879 6556
rect 3879 6500 3883 6556
rect 3819 6496 3883 6500
rect 3899 6556 3963 6560
rect 3899 6500 3903 6556
rect 3903 6500 3959 6556
rect 3959 6500 3963 6556
rect 3899 6496 3963 6500
rect 3979 6556 4043 6560
rect 3979 6500 3983 6556
rect 3983 6500 4039 6556
rect 4039 6500 4043 6556
rect 3979 6496 4043 6500
rect 7994 6556 8058 6560
rect 7994 6500 7998 6556
rect 7998 6500 8054 6556
rect 8054 6500 8058 6556
rect 7994 6496 8058 6500
rect 8074 6556 8138 6560
rect 8074 6500 8078 6556
rect 8078 6500 8134 6556
rect 8134 6500 8138 6556
rect 8074 6496 8138 6500
rect 8154 6556 8218 6560
rect 8154 6500 8158 6556
rect 8158 6500 8214 6556
rect 8214 6500 8218 6556
rect 8154 6496 8218 6500
rect 8234 6556 8298 6560
rect 8234 6500 8238 6556
rect 8238 6500 8294 6556
rect 8294 6500 8298 6556
rect 8234 6496 8298 6500
rect 12249 6556 12313 6560
rect 12249 6500 12253 6556
rect 12253 6500 12309 6556
rect 12309 6500 12313 6556
rect 12249 6496 12313 6500
rect 12329 6556 12393 6560
rect 12329 6500 12333 6556
rect 12333 6500 12389 6556
rect 12389 6500 12393 6556
rect 12329 6496 12393 6500
rect 12409 6556 12473 6560
rect 12409 6500 12413 6556
rect 12413 6500 12469 6556
rect 12469 6500 12473 6556
rect 12409 6496 12473 6500
rect 12489 6556 12553 6560
rect 12489 6500 12493 6556
rect 12493 6500 12549 6556
rect 12549 6500 12553 6556
rect 12489 6496 12553 6500
rect 16504 6556 16568 6560
rect 16504 6500 16508 6556
rect 16508 6500 16564 6556
rect 16564 6500 16568 6556
rect 16504 6496 16568 6500
rect 16584 6556 16648 6560
rect 16584 6500 16588 6556
rect 16588 6500 16644 6556
rect 16644 6500 16648 6556
rect 16584 6496 16648 6500
rect 16664 6556 16728 6560
rect 16664 6500 16668 6556
rect 16668 6500 16724 6556
rect 16724 6500 16728 6556
rect 16664 6496 16728 6500
rect 16744 6556 16808 6560
rect 16744 6500 16748 6556
rect 16748 6500 16804 6556
rect 16804 6500 16808 6556
rect 16744 6496 16808 6500
rect 3079 6012 3143 6016
rect 3079 5956 3083 6012
rect 3083 5956 3139 6012
rect 3139 5956 3143 6012
rect 3079 5952 3143 5956
rect 3159 6012 3223 6016
rect 3159 5956 3163 6012
rect 3163 5956 3219 6012
rect 3219 5956 3223 6012
rect 3159 5952 3223 5956
rect 3239 6012 3303 6016
rect 3239 5956 3243 6012
rect 3243 5956 3299 6012
rect 3299 5956 3303 6012
rect 3239 5952 3303 5956
rect 3319 6012 3383 6016
rect 3319 5956 3323 6012
rect 3323 5956 3379 6012
rect 3379 5956 3383 6012
rect 3319 5952 3383 5956
rect 7334 6012 7398 6016
rect 7334 5956 7338 6012
rect 7338 5956 7394 6012
rect 7394 5956 7398 6012
rect 7334 5952 7398 5956
rect 7414 6012 7478 6016
rect 7414 5956 7418 6012
rect 7418 5956 7474 6012
rect 7474 5956 7478 6012
rect 7414 5952 7478 5956
rect 7494 6012 7558 6016
rect 7494 5956 7498 6012
rect 7498 5956 7554 6012
rect 7554 5956 7558 6012
rect 7494 5952 7558 5956
rect 7574 6012 7638 6016
rect 7574 5956 7578 6012
rect 7578 5956 7634 6012
rect 7634 5956 7638 6012
rect 7574 5952 7638 5956
rect 11589 6012 11653 6016
rect 11589 5956 11593 6012
rect 11593 5956 11649 6012
rect 11649 5956 11653 6012
rect 11589 5952 11653 5956
rect 11669 6012 11733 6016
rect 11669 5956 11673 6012
rect 11673 5956 11729 6012
rect 11729 5956 11733 6012
rect 11669 5952 11733 5956
rect 11749 6012 11813 6016
rect 11749 5956 11753 6012
rect 11753 5956 11809 6012
rect 11809 5956 11813 6012
rect 11749 5952 11813 5956
rect 11829 6012 11893 6016
rect 11829 5956 11833 6012
rect 11833 5956 11889 6012
rect 11889 5956 11893 6012
rect 11829 5952 11893 5956
rect 15844 6012 15908 6016
rect 15844 5956 15848 6012
rect 15848 5956 15904 6012
rect 15904 5956 15908 6012
rect 15844 5952 15908 5956
rect 15924 6012 15988 6016
rect 15924 5956 15928 6012
rect 15928 5956 15984 6012
rect 15984 5956 15988 6012
rect 15924 5952 15988 5956
rect 16004 6012 16068 6016
rect 16004 5956 16008 6012
rect 16008 5956 16064 6012
rect 16064 5956 16068 6012
rect 16004 5952 16068 5956
rect 16084 6012 16148 6016
rect 16084 5956 16088 6012
rect 16088 5956 16144 6012
rect 16144 5956 16148 6012
rect 16084 5952 16148 5956
rect 14412 5808 14476 5812
rect 14412 5752 14426 5808
rect 14426 5752 14476 5808
rect 14412 5748 14476 5752
rect 3739 5468 3803 5472
rect 3739 5412 3743 5468
rect 3743 5412 3799 5468
rect 3799 5412 3803 5468
rect 3739 5408 3803 5412
rect 3819 5468 3883 5472
rect 3819 5412 3823 5468
rect 3823 5412 3879 5468
rect 3879 5412 3883 5468
rect 3819 5408 3883 5412
rect 3899 5468 3963 5472
rect 3899 5412 3903 5468
rect 3903 5412 3959 5468
rect 3959 5412 3963 5468
rect 3899 5408 3963 5412
rect 3979 5468 4043 5472
rect 3979 5412 3983 5468
rect 3983 5412 4039 5468
rect 4039 5412 4043 5468
rect 3979 5408 4043 5412
rect 7994 5468 8058 5472
rect 7994 5412 7998 5468
rect 7998 5412 8054 5468
rect 8054 5412 8058 5468
rect 7994 5408 8058 5412
rect 8074 5468 8138 5472
rect 8074 5412 8078 5468
rect 8078 5412 8134 5468
rect 8134 5412 8138 5468
rect 8074 5408 8138 5412
rect 8154 5468 8218 5472
rect 8154 5412 8158 5468
rect 8158 5412 8214 5468
rect 8214 5412 8218 5468
rect 8154 5408 8218 5412
rect 8234 5468 8298 5472
rect 8234 5412 8238 5468
rect 8238 5412 8294 5468
rect 8294 5412 8298 5468
rect 8234 5408 8298 5412
rect 12249 5468 12313 5472
rect 12249 5412 12253 5468
rect 12253 5412 12309 5468
rect 12309 5412 12313 5468
rect 12249 5408 12313 5412
rect 12329 5468 12393 5472
rect 12329 5412 12333 5468
rect 12333 5412 12389 5468
rect 12389 5412 12393 5468
rect 12329 5408 12393 5412
rect 12409 5468 12473 5472
rect 12409 5412 12413 5468
rect 12413 5412 12469 5468
rect 12469 5412 12473 5468
rect 12409 5408 12473 5412
rect 12489 5468 12553 5472
rect 12489 5412 12493 5468
rect 12493 5412 12549 5468
rect 12549 5412 12553 5468
rect 12489 5408 12553 5412
rect 16504 5468 16568 5472
rect 16504 5412 16508 5468
rect 16508 5412 16564 5468
rect 16564 5412 16568 5468
rect 16504 5408 16568 5412
rect 16584 5468 16648 5472
rect 16584 5412 16588 5468
rect 16588 5412 16644 5468
rect 16644 5412 16648 5468
rect 16584 5408 16648 5412
rect 16664 5468 16728 5472
rect 16664 5412 16668 5468
rect 16668 5412 16724 5468
rect 16724 5412 16728 5468
rect 16664 5408 16728 5412
rect 16744 5468 16808 5472
rect 16744 5412 16748 5468
rect 16748 5412 16804 5468
rect 16804 5412 16808 5468
rect 16744 5408 16808 5412
rect 3079 4924 3143 4928
rect 3079 4868 3083 4924
rect 3083 4868 3139 4924
rect 3139 4868 3143 4924
rect 3079 4864 3143 4868
rect 3159 4924 3223 4928
rect 3159 4868 3163 4924
rect 3163 4868 3219 4924
rect 3219 4868 3223 4924
rect 3159 4864 3223 4868
rect 3239 4924 3303 4928
rect 3239 4868 3243 4924
rect 3243 4868 3299 4924
rect 3299 4868 3303 4924
rect 3239 4864 3303 4868
rect 3319 4924 3383 4928
rect 3319 4868 3323 4924
rect 3323 4868 3379 4924
rect 3379 4868 3383 4924
rect 3319 4864 3383 4868
rect 7334 4924 7398 4928
rect 7334 4868 7338 4924
rect 7338 4868 7394 4924
rect 7394 4868 7398 4924
rect 7334 4864 7398 4868
rect 7414 4924 7478 4928
rect 7414 4868 7418 4924
rect 7418 4868 7474 4924
rect 7474 4868 7478 4924
rect 7414 4864 7478 4868
rect 7494 4924 7558 4928
rect 7494 4868 7498 4924
rect 7498 4868 7554 4924
rect 7554 4868 7558 4924
rect 7494 4864 7558 4868
rect 7574 4924 7638 4928
rect 7574 4868 7578 4924
rect 7578 4868 7634 4924
rect 7634 4868 7638 4924
rect 7574 4864 7638 4868
rect 11589 4924 11653 4928
rect 11589 4868 11593 4924
rect 11593 4868 11649 4924
rect 11649 4868 11653 4924
rect 11589 4864 11653 4868
rect 11669 4924 11733 4928
rect 11669 4868 11673 4924
rect 11673 4868 11729 4924
rect 11729 4868 11733 4924
rect 11669 4864 11733 4868
rect 11749 4924 11813 4928
rect 11749 4868 11753 4924
rect 11753 4868 11809 4924
rect 11809 4868 11813 4924
rect 11749 4864 11813 4868
rect 11829 4924 11893 4928
rect 11829 4868 11833 4924
rect 11833 4868 11889 4924
rect 11889 4868 11893 4924
rect 11829 4864 11893 4868
rect 15844 4924 15908 4928
rect 15844 4868 15848 4924
rect 15848 4868 15904 4924
rect 15904 4868 15908 4924
rect 15844 4864 15908 4868
rect 15924 4924 15988 4928
rect 15924 4868 15928 4924
rect 15928 4868 15984 4924
rect 15984 4868 15988 4924
rect 15924 4864 15988 4868
rect 16004 4924 16068 4928
rect 16004 4868 16008 4924
rect 16008 4868 16064 4924
rect 16064 4868 16068 4924
rect 16004 4864 16068 4868
rect 16084 4924 16148 4928
rect 16084 4868 16088 4924
rect 16088 4868 16144 4924
rect 16144 4868 16148 4924
rect 16084 4864 16148 4868
rect 3739 4380 3803 4384
rect 3739 4324 3743 4380
rect 3743 4324 3799 4380
rect 3799 4324 3803 4380
rect 3739 4320 3803 4324
rect 3819 4380 3883 4384
rect 3819 4324 3823 4380
rect 3823 4324 3879 4380
rect 3879 4324 3883 4380
rect 3819 4320 3883 4324
rect 3899 4380 3963 4384
rect 3899 4324 3903 4380
rect 3903 4324 3959 4380
rect 3959 4324 3963 4380
rect 3899 4320 3963 4324
rect 3979 4380 4043 4384
rect 3979 4324 3983 4380
rect 3983 4324 4039 4380
rect 4039 4324 4043 4380
rect 3979 4320 4043 4324
rect 7994 4380 8058 4384
rect 7994 4324 7998 4380
rect 7998 4324 8054 4380
rect 8054 4324 8058 4380
rect 7994 4320 8058 4324
rect 8074 4380 8138 4384
rect 8074 4324 8078 4380
rect 8078 4324 8134 4380
rect 8134 4324 8138 4380
rect 8074 4320 8138 4324
rect 8154 4380 8218 4384
rect 8154 4324 8158 4380
rect 8158 4324 8214 4380
rect 8214 4324 8218 4380
rect 8154 4320 8218 4324
rect 8234 4380 8298 4384
rect 8234 4324 8238 4380
rect 8238 4324 8294 4380
rect 8294 4324 8298 4380
rect 8234 4320 8298 4324
rect 12249 4380 12313 4384
rect 12249 4324 12253 4380
rect 12253 4324 12309 4380
rect 12309 4324 12313 4380
rect 12249 4320 12313 4324
rect 12329 4380 12393 4384
rect 12329 4324 12333 4380
rect 12333 4324 12389 4380
rect 12389 4324 12393 4380
rect 12329 4320 12393 4324
rect 12409 4380 12473 4384
rect 12409 4324 12413 4380
rect 12413 4324 12469 4380
rect 12469 4324 12473 4380
rect 12409 4320 12473 4324
rect 12489 4380 12553 4384
rect 12489 4324 12493 4380
rect 12493 4324 12549 4380
rect 12549 4324 12553 4380
rect 12489 4320 12553 4324
rect 16504 4380 16568 4384
rect 16504 4324 16508 4380
rect 16508 4324 16564 4380
rect 16564 4324 16568 4380
rect 16504 4320 16568 4324
rect 16584 4380 16648 4384
rect 16584 4324 16588 4380
rect 16588 4324 16644 4380
rect 16644 4324 16648 4380
rect 16584 4320 16648 4324
rect 16664 4380 16728 4384
rect 16664 4324 16668 4380
rect 16668 4324 16724 4380
rect 16724 4324 16728 4380
rect 16664 4320 16728 4324
rect 16744 4380 16808 4384
rect 16744 4324 16748 4380
rect 16748 4324 16804 4380
rect 16804 4324 16808 4380
rect 16744 4320 16808 4324
rect 3079 3836 3143 3840
rect 3079 3780 3083 3836
rect 3083 3780 3139 3836
rect 3139 3780 3143 3836
rect 3079 3776 3143 3780
rect 3159 3836 3223 3840
rect 3159 3780 3163 3836
rect 3163 3780 3219 3836
rect 3219 3780 3223 3836
rect 3159 3776 3223 3780
rect 3239 3836 3303 3840
rect 3239 3780 3243 3836
rect 3243 3780 3299 3836
rect 3299 3780 3303 3836
rect 3239 3776 3303 3780
rect 3319 3836 3383 3840
rect 3319 3780 3323 3836
rect 3323 3780 3379 3836
rect 3379 3780 3383 3836
rect 3319 3776 3383 3780
rect 7334 3836 7398 3840
rect 7334 3780 7338 3836
rect 7338 3780 7394 3836
rect 7394 3780 7398 3836
rect 7334 3776 7398 3780
rect 7414 3836 7478 3840
rect 7414 3780 7418 3836
rect 7418 3780 7474 3836
rect 7474 3780 7478 3836
rect 7414 3776 7478 3780
rect 7494 3836 7558 3840
rect 7494 3780 7498 3836
rect 7498 3780 7554 3836
rect 7554 3780 7558 3836
rect 7494 3776 7558 3780
rect 7574 3836 7638 3840
rect 7574 3780 7578 3836
rect 7578 3780 7634 3836
rect 7634 3780 7638 3836
rect 7574 3776 7638 3780
rect 11589 3836 11653 3840
rect 11589 3780 11593 3836
rect 11593 3780 11649 3836
rect 11649 3780 11653 3836
rect 11589 3776 11653 3780
rect 11669 3836 11733 3840
rect 11669 3780 11673 3836
rect 11673 3780 11729 3836
rect 11729 3780 11733 3836
rect 11669 3776 11733 3780
rect 11749 3836 11813 3840
rect 11749 3780 11753 3836
rect 11753 3780 11809 3836
rect 11809 3780 11813 3836
rect 11749 3776 11813 3780
rect 11829 3836 11893 3840
rect 11829 3780 11833 3836
rect 11833 3780 11889 3836
rect 11889 3780 11893 3836
rect 11829 3776 11893 3780
rect 15844 3836 15908 3840
rect 15844 3780 15848 3836
rect 15848 3780 15904 3836
rect 15904 3780 15908 3836
rect 15844 3776 15908 3780
rect 15924 3836 15988 3840
rect 15924 3780 15928 3836
rect 15928 3780 15984 3836
rect 15984 3780 15988 3836
rect 15924 3776 15988 3780
rect 16004 3836 16068 3840
rect 16004 3780 16008 3836
rect 16008 3780 16064 3836
rect 16064 3780 16068 3836
rect 16004 3776 16068 3780
rect 16084 3836 16148 3840
rect 16084 3780 16088 3836
rect 16088 3780 16144 3836
rect 16144 3780 16148 3836
rect 16084 3776 16148 3780
rect 3739 3292 3803 3296
rect 3739 3236 3743 3292
rect 3743 3236 3799 3292
rect 3799 3236 3803 3292
rect 3739 3232 3803 3236
rect 3819 3292 3883 3296
rect 3819 3236 3823 3292
rect 3823 3236 3879 3292
rect 3879 3236 3883 3292
rect 3819 3232 3883 3236
rect 3899 3292 3963 3296
rect 3899 3236 3903 3292
rect 3903 3236 3959 3292
rect 3959 3236 3963 3292
rect 3899 3232 3963 3236
rect 3979 3292 4043 3296
rect 3979 3236 3983 3292
rect 3983 3236 4039 3292
rect 4039 3236 4043 3292
rect 3979 3232 4043 3236
rect 7994 3292 8058 3296
rect 7994 3236 7998 3292
rect 7998 3236 8054 3292
rect 8054 3236 8058 3292
rect 7994 3232 8058 3236
rect 8074 3292 8138 3296
rect 8074 3236 8078 3292
rect 8078 3236 8134 3292
rect 8134 3236 8138 3292
rect 8074 3232 8138 3236
rect 8154 3292 8218 3296
rect 8154 3236 8158 3292
rect 8158 3236 8214 3292
rect 8214 3236 8218 3292
rect 8154 3232 8218 3236
rect 8234 3292 8298 3296
rect 8234 3236 8238 3292
rect 8238 3236 8294 3292
rect 8294 3236 8298 3292
rect 8234 3232 8298 3236
rect 12249 3292 12313 3296
rect 12249 3236 12253 3292
rect 12253 3236 12309 3292
rect 12309 3236 12313 3292
rect 12249 3232 12313 3236
rect 12329 3292 12393 3296
rect 12329 3236 12333 3292
rect 12333 3236 12389 3292
rect 12389 3236 12393 3292
rect 12329 3232 12393 3236
rect 12409 3292 12473 3296
rect 12409 3236 12413 3292
rect 12413 3236 12469 3292
rect 12469 3236 12473 3292
rect 12409 3232 12473 3236
rect 12489 3292 12553 3296
rect 12489 3236 12493 3292
rect 12493 3236 12549 3292
rect 12549 3236 12553 3292
rect 12489 3232 12553 3236
rect 16504 3292 16568 3296
rect 16504 3236 16508 3292
rect 16508 3236 16564 3292
rect 16564 3236 16568 3292
rect 16504 3232 16568 3236
rect 16584 3292 16648 3296
rect 16584 3236 16588 3292
rect 16588 3236 16644 3292
rect 16644 3236 16648 3292
rect 16584 3232 16648 3236
rect 16664 3292 16728 3296
rect 16664 3236 16668 3292
rect 16668 3236 16724 3292
rect 16724 3236 16728 3292
rect 16664 3232 16728 3236
rect 16744 3292 16808 3296
rect 16744 3236 16748 3292
rect 16748 3236 16804 3292
rect 16804 3236 16808 3292
rect 16744 3232 16808 3236
rect 3079 2748 3143 2752
rect 3079 2692 3083 2748
rect 3083 2692 3139 2748
rect 3139 2692 3143 2748
rect 3079 2688 3143 2692
rect 3159 2748 3223 2752
rect 3159 2692 3163 2748
rect 3163 2692 3219 2748
rect 3219 2692 3223 2748
rect 3159 2688 3223 2692
rect 3239 2748 3303 2752
rect 3239 2692 3243 2748
rect 3243 2692 3299 2748
rect 3299 2692 3303 2748
rect 3239 2688 3303 2692
rect 3319 2748 3383 2752
rect 3319 2692 3323 2748
rect 3323 2692 3379 2748
rect 3379 2692 3383 2748
rect 3319 2688 3383 2692
rect 7334 2748 7398 2752
rect 7334 2692 7338 2748
rect 7338 2692 7394 2748
rect 7394 2692 7398 2748
rect 7334 2688 7398 2692
rect 7414 2748 7478 2752
rect 7414 2692 7418 2748
rect 7418 2692 7474 2748
rect 7474 2692 7478 2748
rect 7414 2688 7478 2692
rect 7494 2748 7558 2752
rect 7494 2692 7498 2748
rect 7498 2692 7554 2748
rect 7554 2692 7558 2748
rect 7494 2688 7558 2692
rect 7574 2748 7638 2752
rect 7574 2692 7578 2748
rect 7578 2692 7634 2748
rect 7634 2692 7638 2748
rect 7574 2688 7638 2692
rect 11589 2748 11653 2752
rect 11589 2692 11593 2748
rect 11593 2692 11649 2748
rect 11649 2692 11653 2748
rect 11589 2688 11653 2692
rect 11669 2748 11733 2752
rect 11669 2692 11673 2748
rect 11673 2692 11729 2748
rect 11729 2692 11733 2748
rect 11669 2688 11733 2692
rect 11749 2748 11813 2752
rect 11749 2692 11753 2748
rect 11753 2692 11809 2748
rect 11809 2692 11813 2748
rect 11749 2688 11813 2692
rect 11829 2748 11893 2752
rect 11829 2692 11833 2748
rect 11833 2692 11889 2748
rect 11889 2692 11893 2748
rect 11829 2688 11893 2692
rect 15844 2748 15908 2752
rect 15844 2692 15848 2748
rect 15848 2692 15904 2748
rect 15904 2692 15908 2748
rect 15844 2688 15908 2692
rect 15924 2748 15988 2752
rect 15924 2692 15928 2748
rect 15928 2692 15984 2748
rect 15984 2692 15988 2748
rect 15924 2688 15988 2692
rect 16004 2748 16068 2752
rect 16004 2692 16008 2748
rect 16008 2692 16064 2748
rect 16064 2692 16068 2748
rect 16004 2688 16068 2692
rect 16084 2748 16148 2752
rect 16084 2692 16088 2748
rect 16088 2692 16144 2748
rect 16144 2692 16148 2748
rect 16084 2688 16148 2692
rect 3739 2204 3803 2208
rect 3739 2148 3743 2204
rect 3743 2148 3799 2204
rect 3799 2148 3803 2204
rect 3739 2144 3803 2148
rect 3819 2204 3883 2208
rect 3819 2148 3823 2204
rect 3823 2148 3879 2204
rect 3879 2148 3883 2204
rect 3819 2144 3883 2148
rect 3899 2204 3963 2208
rect 3899 2148 3903 2204
rect 3903 2148 3959 2204
rect 3959 2148 3963 2204
rect 3899 2144 3963 2148
rect 3979 2204 4043 2208
rect 3979 2148 3983 2204
rect 3983 2148 4039 2204
rect 4039 2148 4043 2204
rect 3979 2144 4043 2148
rect 7994 2204 8058 2208
rect 7994 2148 7998 2204
rect 7998 2148 8054 2204
rect 8054 2148 8058 2204
rect 7994 2144 8058 2148
rect 8074 2204 8138 2208
rect 8074 2148 8078 2204
rect 8078 2148 8134 2204
rect 8134 2148 8138 2204
rect 8074 2144 8138 2148
rect 8154 2204 8218 2208
rect 8154 2148 8158 2204
rect 8158 2148 8214 2204
rect 8214 2148 8218 2204
rect 8154 2144 8218 2148
rect 8234 2204 8298 2208
rect 8234 2148 8238 2204
rect 8238 2148 8294 2204
rect 8294 2148 8298 2204
rect 8234 2144 8298 2148
rect 12249 2204 12313 2208
rect 12249 2148 12253 2204
rect 12253 2148 12309 2204
rect 12309 2148 12313 2204
rect 12249 2144 12313 2148
rect 12329 2204 12393 2208
rect 12329 2148 12333 2204
rect 12333 2148 12389 2204
rect 12389 2148 12393 2204
rect 12329 2144 12393 2148
rect 12409 2204 12473 2208
rect 12409 2148 12413 2204
rect 12413 2148 12469 2204
rect 12469 2148 12473 2204
rect 12409 2144 12473 2148
rect 12489 2204 12553 2208
rect 12489 2148 12493 2204
rect 12493 2148 12549 2204
rect 12549 2148 12553 2204
rect 12489 2144 12553 2148
rect 16504 2204 16568 2208
rect 16504 2148 16508 2204
rect 16508 2148 16564 2204
rect 16564 2148 16568 2204
rect 16504 2144 16568 2148
rect 16584 2204 16648 2208
rect 16584 2148 16588 2204
rect 16588 2148 16644 2204
rect 16644 2148 16648 2204
rect 16584 2144 16648 2148
rect 16664 2204 16728 2208
rect 16664 2148 16668 2204
rect 16668 2148 16724 2204
rect 16724 2148 16728 2204
rect 16664 2144 16728 2148
rect 16744 2204 16808 2208
rect 16744 2148 16748 2204
rect 16748 2148 16804 2204
rect 16804 2148 16808 2204
rect 16744 2144 16808 2148
<< metal4 >>
rect 3071 19072 3391 19088
rect 3071 19008 3079 19072
rect 3143 19008 3159 19072
rect 3223 19008 3239 19072
rect 3303 19008 3319 19072
rect 3383 19008 3391 19072
rect 3071 17984 3391 19008
rect 3071 17920 3079 17984
rect 3143 17920 3159 17984
rect 3223 17920 3239 17984
rect 3303 17920 3319 17984
rect 3383 17920 3391 17984
rect 3071 17050 3391 17920
rect 3731 18528 4051 19088
rect 3731 18464 3739 18528
rect 3803 18464 3819 18528
rect 3883 18464 3899 18528
rect 3963 18464 3979 18528
rect 4043 18464 4051 18528
rect 3555 17780 3621 17781
rect 3555 17716 3556 17780
rect 3620 17716 3621 17780
rect 3555 17715 3621 17716
rect 3071 16896 3113 17050
rect 3349 16896 3391 17050
rect 3071 16832 3079 16896
rect 3383 16832 3391 16896
rect 3071 16814 3113 16832
rect 3349 16814 3391 16832
rect 3071 15808 3391 16814
rect 3071 15744 3079 15808
rect 3143 15744 3159 15808
rect 3223 15744 3239 15808
rect 3303 15744 3319 15808
rect 3383 15744 3391 15808
rect 3071 14720 3391 15744
rect 3071 14656 3079 14720
rect 3143 14656 3159 14720
rect 3223 14656 3239 14720
rect 3303 14656 3319 14720
rect 3383 14656 3391 14720
rect 3071 13632 3391 14656
rect 3071 13568 3079 13632
rect 3143 13568 3159 13632
rect 3223 13568 3239 13632
rect 3303 13568 3319 13632
rect 3383 13568 3391 13632
rect 3071 12834 3391 13568
rect 3071 12598 3113 12834
rect 3349 12598 3391 12834
rect 3071 12544 3391 12598
rect 3071 12480 3079 12544
rect 3143 12480 3159 12544
rect 3223 12480 3239 12544
rect 3303 12480 3319 12544
rect 3383 12480 3391 12544
rect 3071 11456 3391 12480
rect 3071 11392 3079 11456
rect 3143 11392 3159 11456
rect 3223 11392 3239 11456
rect 3303 11392 3319 11456
rect 3383 11392 3391 11456
rect 3071 10368 3391 11392
rect 3558 10709 3618 17715
rect 3731 17710 4051 18464
rect 3731 17474 3773 17710
rect 4009 17474 4051 17710
rect 3731 17440 4051 17474
rect 3731 17376 3739 17440
rect 3803 17376 3819 17440
rect 3883 17376 3899 17440
rect 3963 17376 3979 17440
rect 4043 17376 4051 17440
rect 3731 16352 4051 17376
rect 3731 16288 3739 16352
rect 3803 16288 3819 16352
rect 3883 16288 3899 16352
rect 3963 16288 3979 16352
rect 4043 16288 4051 16352
rect 3731 15264 4051 16288
rect 3731 15200 3739 15264
rect 3803 15200 3819 15264
rect 3883 15200 3899 15264
rect 3963 15200 3979 15264
rect 4043 15200 4051 15264
rect 3731 14176 4051 15200
rect 3731 14112 3739 14176
rect 3803 14112 3819 14176
rect 3883 14112 3899 14176
rect 3963 14112 3979 14176
rect 4043 14112 4051 14176
rect 3731 13494 4051 14112
rect 3731 13258 3773 13494
rect 4009 13258 4051 13494
rect 3731 13088 4051 13258
rect 3731 13024 3739 13088
rect 3803 13024 3819 13088
rect 3883 13024 3899 13088
rect 3963 13024 3979 13088
rect 4043 13024 4051 13088
rect 3731 12000 4051 13024
rect 3731 11936 3739 12000
rect 3803 11936 3819 12000
rect 3883 11936 3899 12000
rect 3963 11936 3979 12000
rect 4043 11936 4051 12000
rect 3731 10912 4051 11936
rect 3731 10848 3739 10912
rect 3803 10848 3819 10912
rect 3883 10848 3899 10912
rect 3963 10848 3979 10912
rect 4043 10848 4051 10912
rect 3555 10708 3621 10709
rect 3555 10644 3556 10708
rect 3620 10644 3621 10708
rect 3555 10643 3621 10644
rect 3071 10304 3079 10368
rect 3143 10304 3159 10368
rect 3223 10304 3239 10368
rect 3303 10304 3319 10368
rect 3383 10304 3391 10368
rect 3071 9280 3391 10304
rect 3071 9216 3079 9280
rect 3143 9216 3159 9280
rect 3223 9216 3239 9280
rect 3303 9216 3319 9280
rect 3383 9216 3391 9280
rect 3071 8618 3391 9216
rect 3071 8382 3113 8618
rect 3349 8382 3391 8618
rect 3071 8192 3391 8382
rect 3071 8128 3079 8192
rect 3143 8128 3159 8192
rect 3223 8128 3239 8192
rect 3303 8128 3319 8192
rect 3383 8128 3391 8192
rect 3071 7104 3391 8128
rect 3071 7040 3079 7104
rect 3143 7040 3159 7104
rect 3223 7040 3239 7104
rect 3303 7040 3319 7104
rect 3383 7040 3391 7104
rect 3071 6016 3391 7040
rect 3071 5952 3079 6016
rect 3143 5952 3159 6016
rect 3223 5952 3239 6016
rect 3303 5952 3319 6016
rect 3383 5952 3391 6016
rect 3071 4928 3391 5952
rect 3071 4864 3079 4928
rect 3143 4864 3159 4928
rect 3223 4864 3239 4928
rect 3303 4864 3319 4928
rect 3383 4864 3391 4928
rect 3071 4402 3391 4864
rect 3071 4166 3113 4402
rect 3349 4166 3391 4402
rect 3071 3840 3391 4166
rect 3071 3776 3079 3840
rect 3143 3776 3159 3840
rect 3223 3776 3239 3840
rect 3303 3776 3319 3840
rect 3383 3776 3391 3840
rect 3071 2752 3391 3776
rect 3071 2688 3079 2752
rect 3143 2688 3159 2752
rect 3223 2688 3239 2752
rect 3303 2688 3319 2752
rect 3383 2688 3391 2752
rect 3071 2128 3391 2688
rect 3731 9824 4051 10848
rect 3731 9760 3739 9824
rect 3803 9760 3819 9824
rect 3883 9760 3899 9824
rect 3963 9760 3979 9824
rect 4043 9760 4051 9824
rect 3731 9278 4051 9760
rect 3731 9042 3773 9278
rect 4009 9042 4051 9278
rect 3731 8736 4051 9042
rect 3731 8672 3739 8736
rect 3803 8672 3819 8736
rect 3883 8672 3899 8736
rect 3963 8672 3979 8736
rect 4043 8672 4051 8736
rect 3731 7648 4051 8672
rect 3731 7584 3739 7648
rect 3803 7584 3819 7648
rect 3883 7584 3899 7648
rect 3963 7584 3979 7648
rect 4043 7584 4051 7648
rect 3731 6560 4051 7584
rect 3731 6496 3739 6560
rect 3803 6496 3819 6560
rect 3883 6496 3899 6560
rect 3963 6496 3979 6560
rect 4043 6496 4051 6560
rect 3731 5472 4051 6496
rect 3731 5408 3739 5472
rect 3803 5408 3819 5472
rect 3883 5408 3899 5472
rect 3963 5408 3979 5472
rect 4043 5408 4051 5472
rect 3731 5062 4051 5408
rect 3731 4826 3773 5062
rect 4009 4826 4051 5062
rect 3731 4384 4051 4826
rect 3731 4320 3739 4384
rect 3803 4320 3819 4384
rect 3883 4320 3899 4384
rect 3963 4320 3979 4384
rect 4043 4320 4051 4384
rect 3731 3296 4051 4320
rect 3731 3232 3739 3296
rect 3803 3232 3819 3296
rect 3883 3232 3899 3296
rect 3963 3232 3979 3296
rect 4043 3232 4051 3296
rect 3731 2208 4051 3232
rect 3731 2144 3739 2208
rect 3803 2144 3819 2208
rect 3883 2144 3899 2208
rect 3963 2144 3979 2208
rect 4043 2144 4051 2208
rect 3731 2128 4051 2144
rect 7326 19072 7646 19088
rect 7326 19008 7334 19072
rect 7398 19008 7414 19072
rect 7478 19008 7494 19072
rect 7558 19008 7574 19072
rect 7638 19008 7646 19072
rect 7326 17984 7646 19008
rect 7326 17920 7334 17984
rect 7398 17920 7414 17984
rect 7478 17920 7494 17984
rect 7558 17920 7574 17984
rect 7638 17920 7646 17984
rect 7326 17050 7646 17920
rect 7326 16896 7368 17050
rect 7604 16896 7646 17050
rect 7326 16832 7334 16896
rect 7638 16832 7646 16896
rect 7326 16814 7368 16832
rect 7604 16814 7646 16832
rect 7326 15808 7646 16814
rect 7326 15744 7334 15808
rect 7398 15744 7414 15808
rect 7478 15744 7494 15808
rect 7558 15744 7574 15808
rect 7638 15744 7646 15808
rect 7326 14720 7646 15744
rect 7326 14656 7334 14720
rect 7398 14656 7414 14720
rect 7478 14656 7494 14720
rect 7558 14656 7574 14720
rect 7638 14656 7646 14720
rect 7326 13632 7646 14656
rect 7326 13568 7334 13632
rect 7398 13568 7414 13632
rect 7478 13568 7494 13632
rect 7558 13568 7574 13632
rect 7638 13568 7646 13632
rect 7326 12834 7646 13568
rect 7326 12598 7368 12834
rect 7604 12598 7646 12834
rect 7326 12544 7646 12598
rect 7326 12480 7334 12544
rect 7398 12480 7414 12544
rect 7478 12480 7494 12544
rect 7558 12480 7574 12544
rect 7638 12480 7646 12544
rect 7326 11456 7646 12480
rect 7326 11392 7334 11456
rect 7398 11392 7414 11456
rect 7478 11392 7494 11456
rect 7558 11392 7574 11456
rect 7638 11392 7646 11456
rect 7326 10368 7646 11392
rect 7326 10304 7334 10368
rect 7398 10304 7414 10368
rect 7478 10304 7494 10368
rect 7558 10304 7574 10368
rect 7638 10304 7646 10368
rect 7326 9280 7646 10304
rect 7326 9216 7334 9280
rect 7398 9216 7414 9280
rect 7478 9216 7494 9280
rect 7558 9216 7574 9280
rect 7638 9216 7646 9280
rect 7326 8618 7646 9216
rect 7326 8382 7368 8618
rect 7604 8382 7646 8618
rect 7326 8192 7646 8382
rect 7326 8128 7334 8192
rect 7398 8128 7414 8192
rect 7478 8128 7494 8192
rect 7558 8128 7574 8192
rect 7638 8128 7646 8192
rect 7326 7104 7646 8128
rect 7326 7040 7334 7104
rect 7398 7040 7414 7104
rect 7478 7040 7494 7104
rect 7558 7040 7574 7104
rect 7638 7040 7646 7104
rect 7326 6016 7646 7040
rect 7326 5952 7334 6016
rect 7398 5952 7414 6016
rect 7478 5952 7494 6016
rect 7558 5952 7574 6016
rect 7638 5952 7646 6016
rect 7326 4928 7646 5952
rect 7326 4864 7334 4928
rect 7398 4864 7414 4928
rect 7478 4864 7494 4928
rect 7558 4864 7574 4928
rect 7638 4864 7646 4928
rect 7326 4402 7646 4864
rect 7326 4166 7368 4402
rect 7604 4166 7646 4402
rect 7326 3840 7646 4166
rect 7326 3776 7334 3840
rect 7398 3776 7414 3840
rect 7478 3776 7494 3840
rect 7558 3776 7574 3840
rect 7638 3776 7646 3840
rect 7326 2752 7646 3776
rect 7326 2688 7334 2752
rect 7398 2688 7414 2752
rect 7478 2688 7494 2752
rect 7558 2688 7574 2752
rect 7638 2688 7646 2752
rect 7326 2128 7646 2688
rect 7986 18528 8306 19088
rect 7986 18464 7994 18528
rect 8058 18464 8074 18528
rect 8138 18464 8154 18528
rect 8218 18464 8234 18528
rect 8298 18464 8306 18528
rect 7986 17710 8306 18464
rect 7986 17474 8028 17710
rect 8264 17474 8306 17710
rect 7986 17440 8306 17474
rect 7986 17376 7994 17440
rect 8058 17376 8074 17440
rect 8138 17376 8154 17440
rect 8218 17376 8234 17440
rect 8298 17376 8306 17440
rect 7986 16352 8306 17376
rect 7986 16288 7994 16352
rect 8058 16288 8074 16352
rect 8138 16288 8154 16352
rect 8218 16288 8234 16352
rect 8298 16288 8306 16352
rect 7986 15264 8306 16288
rect 7986 15200 7994 15264
rect 8058 15200 8074 15264
rect 8138 15200 8154 15264
rect 8218 15200 8234 15264
rect 8298 15200 8306 15264
rect 7986 14176 8306 15200
rect 7986 14112 7994 14176
rect 8058 14112 8074 14176
rect 8138 14112 8154 14176
rect 8218 14112 8234 14176
rect 8298 14112 8306 14176
rect 7986 13494 8306 14112
rect 11581 19072 11901 19088
rect 11581 19008 11589 19072
rect 11653 19008 11669 19072
rect 11733 19008 11749 19072
rect 11813 19008 11829 19072
rect 11893 19008 11901 19072
rect 11581 17984 11901 19008
rect 11581 17920 11589 17984
rect 11653 17920 11669 17984
rect 11733 17920 11749 17984
rect 11813 17920 11829 17984
rect 11893 17920 11901 17984
rect 11581 17050 11901 17920
rect 11581 16896 11623 17050
rect 11859 16896 11901 17050
rect 11581 16832 11589 16896
rect 11893 16832 11901 16896
rect 11581 16814 11623 16832
rect 11859 16814 11901 16832
rect 11581 15808 11901 16814
rect 11581 15744 11589 15808
rect 11653 15744 11669 15808
rect 11733 15744 11749 15808
rect 11813 15744 11829 15808
rect 11893 15744 11901 15808
rect 11581 14720 11901 15744
rect 11581 14656 11589 14720
rect 11653 14656 11669 14720
rect 11733 14656 11749 14720
rect 11813 14656 11829 14720
rect 11893 14656 11901 14720
rect 10731 13836 10797 13837
rect 10731 13772 10732 13836
rect 10796 13772 10797 13836
rect 10731 13771 10797 13772
rect 7986 13258 8028 13494
rect 8264 13258 8306 13494
rect 10734 13429 10794 13771
rect 11581 13632 11901 14656
rect 11581 13568 11589 13632
rect 11653 13568 11669 13632
rect 11733 13568 11749 13632
rect 11813 13568 11829 13632
rect 11893 13568 11901 13632
rect 10731 13428 10797 13429
rect 10731 13364 10732 13428
rect 10796 13364 10797 13428
rect 10731 13363 10797 13364
rect 7986 13088 8306 13258
rect 7986 13024 7994 13088
rect 8058 13024 8074 13088
rect 8138 13024 8154 13088
rect 8218 13024 8234 13088
rect 8298 13024 8306 13088
rect 7986 12000 8306 13024
rect 7986 11936 7994 12000
rect 8058 11936 8074 12000
rect 8138 11936 8154 12000
rect 8218 11936 8234 12000
rect 8298 11936 8306 12000
rect 7986 10912 8306 11936
rect 7986 10848 7994 10912
rect 8058 10848 8074 10912
rect 8138 10848 8154 10912
rect 8218 10848 8234 10912
rect 8298 10848 8306 10912
rect 7986 9824 8306 10848
rect 10734 10845 10794 13363
rect 11581 12834 11901 13568
rect 11581 12598 11623 12834
rect 11859 12598 11901 12834
rect 11581 12544 11901 12598
rect 11581 12480 11589 12544
rect 11653 12480 11669 12544
rect 11733 12480 11749 12544
rect 11813 12480 11829 12544
rect 11893 12480 11901 12544
rect 11581 11456 11901 12480
rect 11581 11392 11589 11456
rect 11653 11392 11669 11456
rect 11733 11392 11749 11456
rect 11813 11392 11829 11456
rect 11893 11392 11901 11456
rect 10731 10844 10797 10845
rect 10731 10780 10732 10844
rect 10796 10780 10797 10844
rect 10731 10779 10797 10780
rect 7986 9760 7994 9824
rect 8058 9760 8074 9824
rect 8138 9760 8154 9824
rect 8218 9760 8234 9824
rect 8298 9760 8306 9824
rect 7986 9278 8306 9760
rect 7986 9042 8028 9278
rect 8264 9042 8306 9278
rect 7986 8736 8306 9042
rect 7986 8672 7994 8736
rect 8058 8672 8074 8736
rect 8138 8672 8154 8736
rect 8218 8672 8234 8736
rect 8298 8672 8306 8736
rect 7986 7648 8306 8672
rect 10734 7989 10794 10779
rect 11581 10368 11901 11392
rect 11581 10304 11589 10368
rect 11653 10304 11669 10368
rect 11733 10304 11749 10368
rect 11813 10304 11829 10368
rect 11893 10304 11901 10368
rect 11581 9280 11901 10304
rect 11581 9216 11589 9280
rect 11653 9216 11669 9280
rect 11733 9216 11749 9280
rect 11813 9216 11829 9280
rect 11893 9216 11901 9280
rect 11581 8618 11901 9216
rect 11581 8382 11623 8618
rect 11859 8382 11901 8618
rect 11581 8192 11901 8382
rect 11581 8128 11589 8192
rect 11653 8128 11669 8192
rect 11733 8128 11749 8192
rect 11813 8128 11829 8192
rect 11893 8128 11901 8192
rect 10731 7988 10797 7989
rect 10731 7924 10732 7988
rect 10796 7924 10797 7988
rect 10731 7923 10797 7924
rect 7986 7584 7994 7648
rect 8058 7584 8074 7648
rect 8138 7584 8154 7648
rect 8218 7584 8234 7648
rect 8298 7584 8306 7648
rect 7986 6560 8306 7584
rect 7986 6496 7994 6560
rect 8058 6496 8074 6560
rect 8138 6496 8154 6560
rect 8218 6496 8234 6560
rect 8298 6496 8306 6560
rect 7986 5472 8306 6496
rect 7986 5408 7994 5472
rect 8058 5408 8074 5472
rect 8138 5408 8154 5472
rect 8218 5408 8234 5472
rect 8298 5408 8306 5472
rect 7986 5062 8306 5408
rect 7986 4826 8028 5062
rect 8264 4826 8306 5062
rect 7986 4384 8306 4826
rect 7986 4320 7994 4384
rect 8058 4320 8074 4384
rect 8138 4320 8154 4384
rect 8218 4320 8234 4384
rect 8298 4320 8306 4384
rect 7986 3296 8306 4320
rect 7986 3232 7994 3296
rect 8058 3232 8074 3296
rect 8138 3232 8154 3296
rect 8218 3232 8234 3296
rect 8298 3232 8306 3296
rect 7986 2208 8306 3232
rect 7986 2144 7994 2208
rect 8058 2144 8074 2208
rect 8138 2144 8154 2208
rect 8218 2144 8234 2208
rect 8298 2144 8306 2208
rect 7986 2128 8306 2144
rect 11581 7104 11901 8128
rect 11581 7040 11589 7104
rect 11653 7040 11669 7104
rect 11733 7040 11749 7104
rect 11813 7040 11829 7104
rect 11893 7040 11901 7104
rect 11581 6016 11901 7040
rect 11581 5952 11589 6016
rect 11653 5952 11669 6016
rect 11733 5952 11749 6016
rect 11813 5952 11829 6016
rect 11893 5952 11901 6016
rect 11581 4928 11901 5952
rect 11581 4864 11589 4928
rect 11653 4864 11669 4928
rect 11733 4864 11749 4928
rect 11813 4864 11829 4928
rect 11893 4864 11901 4928
rect 11581 4402 11901 4864
rect 11581 4166 11623 4402
rect 11859 4166 11901 4402
rect 11581 3840 11901 4166
rect 11581 3776 11589 3840
rect 11653 3776 11669 3840
rect 11733 3776 11749 3840
rect 11813 3776 11829 3840
rect 11893 3776 11901 3840
rect 11581 2752 11901 3776
rect 11581 2688 11589 2752
rect 11653 2688 11669 2752
rect 11733 2688 11749 2752
rect 11813 2688 11829 2752
rect 11893 2688 11901 2752
rect 11581 2128 11901 2688
rect 12241 18528 12561 19088
rect 12241 18464 12249 18528
rect 12313 18464 12329 18528
rect 12393 18464 12409 18528
rect 12473 18464 12489 18528
rect 12553 18464 12561 18528
rect 12241 17710 12561 18464
rect 12241 17474 12283 17710
rect 12519 17474 12561 17710
rect 12241 17440 12561 17474
rect 12241 17376 12249 17440
rect 12313 17376 12329 17440
rect 12393 17376 12409 17440
rect 12473 17376 12489 17440
rect 12553 17376 12561 17440
rect 12241 16352 12561 17376
rect 12241 16288 12249 16352
rect 12313 16288 12329 16352
rect 12393 16288 12409 16352
rect 12473 16288 12489 16352
rect 12553 16288 12561 16352
rect 12241 15264 12561 16288
rect 12241 15200 12249 15264
rect 12313 15200 12329 15264
rect 12393 15200 12409 15264
rect 12473 15200 12489 15264
rect 12553 15200 12561 15264
rect 12241 14176 12561 15200
rect 15836 19072 16156 19088
rect 15836 19008 15844 19072
rect 15908 19008 15924 19072
rect 15988 19008 16004 19072
rect 16068 19008 16084 19072
rect 16148 19008 16156 19072
rect 15836 17984 16156 19008
rect 15836 17920 15844 17984
rect 15908 17920 15924 17984
rect 15988 17920 16004 17984
rect 16068 17920 16084 17984
rect 16148 17920 16156 17984
rect 15836 17050 16156 17920
rect 15836 16896 15878 17050
rect 16114 16896 16156 17050
rect 15836 16832 15844 16896
rect 16148 16832 16156 16896
rect 15836 16814 15878 16832
rect 16114 16814 16156 16832
rect 15836 15808 16156 16814
rect 15836 15744 15844 15808
rect 15908 15744 15924 15808
rect 15988 15744 16004 15808
rect 16068 15744 16084 15808
rect 16148 15744 16156 15808
rect 12755 15060 12821 15061
rect 12755 14996 12756 15060
rect 12820 14996 12821 15060
rect 12755 14995 12821 14996
rect 12241 14112 12249 14176
rect 12313 14112 12329 14176
rect 12393 14112 12409 14176
rect 12473 14112 12489 14176
rect 12553 14112 12561 14176
rect 12241 13494 12561 14112
rect 12241 13258 12283 13494
rect 12519 13258 12561 13494
rect 12241 13088 12561 13258
rect 12241 13024 12249 13088
rect 12313 13024 12329 13088
rect 12393 13024 12409 13088
rect 12473 13024 12489 13088
rect 12553 13024 12561 13088
rect 12241 12000 12561 13024
rect 12241 11936 12249 12000
rect 12313 11936 12329 12000
rect 12393 11936 12409 12000
rect 12473 11936 12489 12000
rect 12553 11936 12561 12000
rect 12241 10912 12561 11936
rect 12241 10848 12249 10912
rect 12313 10848 12329 10912
rect 12393 10848 12409 10912
rect 12473 10848 12489 10912
rect 12553 10848 12561 10912
rect 12241 9824 12561 10848
rect 12758 10301 12818 14995
rect 14411 14788 14477 14789
rect 14411 14724 14412 14788
rect 14476 14724 14477 14788
rect 14411 14723 14477 14724
rect 12755 10300 12821 10301
rect 12755 10236 12756 10300
rect 12820 10236 12821 10300
rect 12755 10235 12821 10236
rect 12241 9760 12249 9824
rect 12313 9760 12329 9824
rect 12393 9760 12409 9824
rect 12473 9760 12489 9824
rect 12553 9760 12561 9824
rect 12241 9278 12561 9760
rect 12241 9042 12283 9278
rect 12519 9042 12561 9278
rect 12241 8736 12561 9042
rect 12241 8672 12249 8736
rect 12313 8672 12329 8736
rect 12393 8672 12409 8736
rect 12473 8672 12489 8736
rect 12553 8672 12561 8736
rect 12241 7648 12561 8672
rect 12241 7584 12249 7648
rect 12313 7584 12329 7648
rect 12393 7584 12409 7648
rect 12473 7584 12489 7648
rect 12553 7584 12561 7648
rect 12241 6560 12561 7584
rect 12241 6496 12249 6560
rect 12313 6496 12329 6560
rect 12393 6496 12409 6560
rect 12473 6496 12489 6560
rect 12553 6496 12561 6560
rect 12241 5472 12561 6496
rect 14414 5813 14474 14723
rect 15836 14720 16156 15744
rect 15836 14656 15844 14720
rect 15908 14656 15924 14720
rect 15988 14656 16004 14720
rect 16068 14656 16084 14720
rect 16148 14656 16156 14720
rect 15836 13632 16156 14656
rect 15836 13568 15844 13632
rect 15908 13568 15924 13632
rect 15988 13568 16004 13632
rect 16068 13568 16084 13632
rect 16148 13568 16156 13632
rect 15836 12834 16156 13568
rect 15836 12598 15878 12834
rect 16114 12598 16156 12834
rect 15836 12544 16156 12598
rect 15836 12480 15844 12544
rect 15908 12480 15924 12544
rect 15988 12480 16004 12544
rect 16068 12480 16084 12544
rect 16148 12480 16156 12544
rect 15836 11456 16156 12480
rect 15836 11392 15844 11456
rect 15908 11392 15924 11456
rect 15988 11392 16004 11456
rect 16068 11392 16084 11456
rect 16148 11392 16156 11456
rect 15836 10368 16156 11392
rect 15836 10304 15844 10368
rect 15908 10304 15924 10368
rect 15988 10304 16004 10368
rect 16068 10304 16084 10368
rect 16148 10304 16156 10368
rect 15836 9280 16156 10304
rect 15836 9216 15844 9280
rect 15908 9216 15924 9280
rect 15988 9216 16004 9280
rect 16068 9216 16084 9280
rect 16148 9216 16156 9280
rect 15836 8618 16156 9216
rect 15836 8382 15878 8618
rect 16114 8382 16156 8618
rect 15836 8192 16156 8382
rect 15836 8128 15844 8192
rect 15908 8128 15924 8192
rect 15988 8128 16004 8192
rect 16068 8128 16084 8192
rect 16148 8128 16156 8192
rect 15836 7104 16156 8128
rect 15836 7040 15844 7104
rect 15908 7040 15924 7104
rect 15988 7040 16004 7104
rect 16068 7040 16084 7104
rect 16148 7040 16156 7104
rect 15836 6016 16156 7040
rect 15836 5952 15844 6016
rect 15908 5952 15924 6016
rect 15988 5952 16004 6016
rect 16068 5952 16084 6016
rect 16148 5952 16156 6016
rect 14411 5812 14477 5813
rect 14411 5748 14412 5812
rect 14476 5748 14477 5812
rect 14411 5747 14477 5748
rect 12241 5408 12249 5472
rect 12313 5408 12329 5472
rect 12393 5408 12409 5472
rect 12473 5408 12489 5472
rect 12553 5408 12561 5472
rect 12241 5062 12561 5408
rect 12241 4826 12283 5062
rect 12519 4826 12561 5062
rect 12241 4384 12561 4826
rect 12241 4320 12249 4384
rect 12313 4320 12329 4384
rect 12393 4320 12409 4384
rect 12473 4320 12489 4384
rect 12553 4320 12561 4384
rect 12241 3296 12561 4320
rect 12241 3232 12249 3296
rect 12313 3232 12329 3296
rect 12393 3232 12409 3296
rect 12473 3232 12489 3296
rect 12553 3232 12561 3296
rect 12241 2208 12561 3232
rect 12241 2144 12249 2208
rect 12313 2144 12329 2208
rect 12393 2144 12409 2208
rect 12473 2144 12489 2208
rect 12553 2144 12561 2208
rect 12241 2128 12561 2144
rect 15836 4928 16156 5952
rect 15836 4864 15844 4928
rect 15908 4864 15924 4928
rect 15988 4864 16004 4928
rect 16068 4864 16084 4928
rect 16148 4864 16156 4928
rect 15836 4402 16156 4864
rect 15836 4166 15878 4402
rect 16114 4166 16156 4402
rect 15836 3840 16156 4166
rect 15836 3776 15844 3840
rect 15908 3776 15924 3840
rect 15988 3776 16004 3840
rect 16068 3776 16084 3840
rect 16148 3776 16156 3840
rect 15836 2752 16156 3776
rect 15836 2688 15844 2752
rect 15908 2688 15924 2752
rect 15988 2688 16004 2752
rect 16068 2688 16084 2752
rect 16148 2688 16156 2752
rect 15836 2128 16156 2688
rect 16496 18528 16816 19088
rect 16496 18464 16504 18528
rect 16568 18464 16584 18528
rect 16648 18464 16664 18528
rect 16728 18464 16744 18528
rect 16808 18464 16816 18528
rect 16496 17710 16816 18464
rect 16496 17474 16538 17710
rect 16774 17474 16816 17710
rect 16496 17440 16816 17474
rect 16496 17376 16504 17440
rect 16568 17376 16584 17440
rect 16648 17376 16664 17440
rect 16728 17376 16744 17440
rect 16808 17376 16816 17440
rect 16496 16352 16816 17376
rect 16496 16288 16504 16352
rect 16568 16288 16584 16352
rect 16648 16288 16664 16352
rect 16728 16288 16744 16352
rect 16808 16288 16816 16352
rect 16496 15264 16816 16288
rect 16496 15200 16504 15264
rect 16568 15200 16584 15264
rect 16648 15200 16664 15264
rect 16728 15200 16744 15264
rect 16808 15200 16816 15264
rect 16496 14176 16816 15200
rect 16496 14112 16504 14176
rect 16568 14112 16584 14176
rect 16648 14112 16664 14176
rect 16728 14112 16744 14176
rect 16808 14112 16816 14176
rect 16496 13494 16816 14112
rect 16496 13258 16538 13494
rect 16774 13258 16816 13494
rect 16496 13088 16816 13258
rect 16496 13024 16504 13088
rect 16568 13024 16584 13088
rect 16648 13024 16664 13088
rect 16728 13024 16744 13088
rect 16808 13024 16816 13088
rect 16496 12000 16816 13024
rect 16496 11936 16504 12000
rect 16568 11936 16584 12000
rect 16648 11936 16664 12000
rect 16728 11936 16744 12000
rect 16808 11936 16816 12000
rect 16496 10912 16816 11936
rect 16496 10848 16504 10912
rect 16568 10848 16584 10912
rect 16648 10848 16664 10912
rect 16728 10848 16744 10912
rect 16808 10848 16816 10912
rect 16496 9824 16816 10848
rect 16496 9760 16504 9824
rect 16568 9760 16584 9824
rect 16648 9760 16664 9824
rect 16728 9760 16744 9824
rect 16808 9760 16816 9824
rect 16496 9278 16816 9760
rect 16496 9042 16538 9278
rect 16774 9042 16816 9278
rect 16496 8736 16816 9042
rect 16496 8672 16504 8736
rect 16568 8672 16584 8736
rect 16648 8672 16664 8736
rect 16728 8672 16744 8736
rect 16808 8672 16816 8736
rect 16496 7648 16816 8672
rect 16496 7584 16504 7648
rect 16568 7584 16584 7648
rect 16648 7584 16664 7648
rect 16728 7584 16744 7648
rect 16808 7584 16816 7648
rect 16496 6560 16816 7584
rect 16496 6496 16504 6560
rect 16568 6496 16584 6560
rect 16648 6496 16664 6560
rect 16728 6496 16744 6560
rect 16808 6496 16816 6560
rect 16496 5472 16816 6496
rect 16496 5408 16504 5472
rect 16568 5408 16584 5472
rect 16648 5408 16664 5472
rect 16728 5408 16744 5472
rect 16808 5408 16816 5472
rect 16496 5062 16816 5408
rect 16496 4826 16538 5062
rect 16774 4826 16816 5062
rect 16496 4384 16816 4826
rect 16496 4320 16504 4384
rect 16568 4320 16584 4384
rect 16648 4320 16664 4384
rect 16728 4320 16744 4384
rect 16808 4320 16816 4384
rect 16496 3296 16816 4320
rect 16496 3232 16504 3296
rect 16568 3232 16584 3296
rect 16648 3232 16664 3296
rect 16728 3232 16744 3296
rect 16808 3232 16816 3296
rect 16496 2208 16816 3232
rect 16496 2144 16504 2208
rect 16568 2144 16584 2208
rect 16648 2144 16664 2208
rect 16728 2144 16744 2208
rect 16808 2144 16816 2208
rect 16496 2128 16816 2144
<< via4 >>
rect 3113 16896 3349 17050
rect 3113 16832 3143 16896
rect 3143 16832 3159 16896
rect 3159 16832 3223 16896
rect 3223 16832 3239 16896
rect 3239 16832 3303 16896
rect 3303 16832 3319 16896
rect 3319 16832 3349 16896
rect 3113 16814 3349 16832
rect 3113 12598 3349 12834
rect 3773 17474 4009 17710
rect 3773 13258 4009 13494
rect 3113 8382 3349 8618
rect 3113 4166 3349 4402
rect 3773 9042 4009 9278
rect 3773 4826 4009 5062
rect 7368 16896 7604 17050
rect 7368 16832 7398 16896
rect 7398 16832 7414 16896
rect 7414 16832 7478 16896
rect 7478 16832 7494 16896
rect 7494 16832 7558 16896
rect 7558 16832 7574 16896
rect 7574 16832 7604 16896
rect 7368 16814 7604 16832
rect 7368 12598 7604 12834
rect 7368 8382 7604 8618
rect 7368 4166 7604 4402
rect 8028 17474 8264 17710
rect 11623 16896 11859 17050
rect 11623 16832 11653 16896
rect 11653 16832 11669 16896
rect 11669 16832 11733 16896
rect 11733 16832 11749 16896
rect 11749 16832 11813 16896
rect 11813 16832 11829 16896
rect 11829 16832 11859 16896
rect 11623 16814 11859 16832
rect 8028 13258 8264 13494
rect 11623 12598 11859 12834
rect 8028 9042 8264 9278
rect 11623 8382 11859 8618
rect 8028 4826 8264 5062
rect 11623 4166 11859 4402
rect 12283 17474 12519 17710
rect 15878 16896 16114 17050
rect 15878 16832 15908 16896
rect 15908 16832 15924 16896
rect 15924 16832 15988 16896
rect 15988 16832 16004 16896
rect 16004 16832 16068 16896
rect 16068 16832 16084 16896
rect 16084 16832 16114 16896
rect 15878 16814 16114 16832
rect 12283 13258 12519 13494
rect 12283 9042 12519 9278
rect 15878 12598 16114 12834
rect 15878 8382 16114 8618
rect 12283 4826 12519 5062
rect 15878 4166 16114 4402
rect 16538 17474 16774 17710
rect 16538 13258 16774 13494
rect 16538 9042 16774 9278
rect 16538 4826 16774 5062
<< metal5 >>
rect 1056 17710 18172 17752
rect 1056 17474 3773 17710
rect 4009 17474 8028 17710
rect 8264 17474 12283 17710
rect 12519 17474 16538 17710
rect 16774 17474 18172 17710
rect 1056 17432 18172 17474
rect 1056 17050 18172 17092
rect 1056 16814 3113 17050
rect 3349 16814 7368 17050
rect 7604 16814 11623 17050
rect 11859 16814 15878 17050
rect 16114 16814 18172 17050
rect 1056 16772 18172 16814
rect 1056 13494 18172 13536
rect 1056 13258 3773 13494
rect 4009 13258 8028 13494
rect 8264 13258 12283 13494
rect 12519 13258 16538 13494
rect 16774 13258 18172 13494
rect 1056 13216 18172 13258
rect 1056 12834 18172 12876
rect 1056 12598 3113 12834
rect 3349 12598 7368 12834
rect 7604 12598 11623 12834
rect 11859 12598 15878 12834
rect 16114 12598 18172 12834
rect 1056 12556 18172 12598
rect 1056 9278 18172 9320
rect 1056 9042 3773 9278
rect 4009 9042 8028 9278
rect 8264 9042 12283 9278
rect 12519 9042 16538 9278
rect 16774 9042 18172 9278
rect 1056 9000 18172 9042
rect 1056 8618 18172 8660
rect 1056 8382 3113 8618
rect 3349 8382 7368 8618
rect 7604 8382 11623 8618
rect 11859 8382 15878 8618
rect 16114 8382 18172 8618
rect 1056 8340 18172 8382
rect 1056 5062 18172 5104
rect 1056 4826 3773 5062
rect 4009 4826 8028 5062
rect 8264 4826 12283 5062
rect 12519 4826 16538 5062
rect 16774 4826 18172 5062
rect 1056 4784 18172 4826
rect 1056 4402 18172 4444
rect 1056 4166 3113 4402
rect 3349 4166 7368 4402
rect 7604 4166 11623 4402
rect 11859 4166 15878 4402
rect 16114 4166 18172 4402
rect 1056 4124 18172 4166
use sky130_fd_sc_hd__inv_2  _233_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8372 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _234_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12236 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _235_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12052 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _236_
timestamp 1704896540
transform 1 0 13156 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _237_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _238_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5244 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _239_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 15272 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _240_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _241_
timestamp 1704896540
transform -1 0 15732 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _242_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 3772 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _243_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 7084 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _244_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 6348 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _245_
timestamp 1704896540
transform 1 0 4692 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _246_
timestamp 1704896540
transform 1 0 4968 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _247_
timestamp 1704896540
transform 1 0 6440 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _248_
timestamp 1704896540
transform -1 0 3680 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _249_
timestamp 1704896540
transform 1 0 5612 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _250_
timestamp 1704896540
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _251_
timestamp 1704896540
transform 1 0 6348 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _252_
timestamp 1704896540
transform -1 0 7636 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _253_
timestamp 1704896540
transform 1 0 6624 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _254_
timestamp 1704896540
transform -1 0 4600 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _255_
timestamp 1704896540
transform 1 0 5888 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _256_
timestamp 1704896540
transform 1 0 6624 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _257_
timestamp 1704896540
transform 1 0 8556 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _258_
timestamp 1704896540
transform 1 0 9200 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _259_
timestamp 1704896540
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _260_
timestamp 1704896540
transform 1 0 9660 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _261_
timestamp 1704896540
transform 1 0 9752 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _262_
timestamp 1704896540
transform 1 0 9936 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _263_
timestamp 1704896540
transform -1 0 16008 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _264_
timestamp 1704896540
transform 1 0 12788 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _265_
timestamp 1704896540
transform 1 0 14076 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _266_
timestamp 1704896540
transform 1 0 15548 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _267_
timestamp 1704896540
transform 1 0 13984 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _268_
timestamp 1704896540
transform -1 0 14720 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _269_
timestamp 1704896540
transform 1 0 11868 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _270_
timestamp 1704896540
transform 1 0 12604 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _271_
timestamp 1704896540
transform -1 0 13984 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _272_
timestamp 1704896540
transform 1 0 14720 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _273_
timestamp 1704896540
transform -1 0 14536 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _274_
timestamp 1704896540
transform -1 0 13708 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _275_
timestamp 1704896540
transform 1 0 12788 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _276_
timestamp 1704896540
transform -1 0 14628 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _277_
timestamp 1704896540
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _278_
timestamp 1704896540
transform 1 0 14076 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _279_
timestamp 1704896540
transform 1 0 12328 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _280_
timestamp 1704896540
transform -1 0 13984 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _281_
timestamp 1704896540
transform 1 0 9200 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _282_
timestamp 1704896540
transform 1 0 9936 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _283_
timestamp 1704896540
transform 1 0 11224 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _284_
timestamp 1704896540
transform 1 0 11592 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _285_
timestamp 1704896540
transform 1 0 10488 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _286_
timestamp 1704896540
transform -1 0 11224 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1704896540
transform 1 0 8924 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _288_
timestamp 1704896540
transform -1 0 14628 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _289_
timestamp 1704896540
transform 1 0 12604 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _290_
timestamp 1704896540
transform 1 0 12880 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _291_
timestamp 1704896540
transform 1 0 4324 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _292_
timestamp 1704896540
transform -1 0 6348 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _293_
timestamp 1704896540
transform -1 0 12604 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__o21ba_1  _294_
timestamp 1704896540
transform 1 0 6348 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _295_
timestamp 1704896540
transform -1 0 15180 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _296_
timestamp 1704896540
transform -1 0 3680 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _297_
timestamp 1704896540
transform 1 0 5520 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _298_
timestamp 1704896540
transform 1 0 6072 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _299_
timestamp 1704896540
transform 1 0 4324 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _300_
timestamp 1704896540
transform 1 0 5060 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _301_
timestamp 1704896540
transform 1 0 6348 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _302_
timestamp 1704896540
transform -1 0 4140 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _303_
timestamp 1704896540
transform 1 0 5520 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _304_
timestamp 1704896540
transform 1 0 7728 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _305_
timestamp 1704896540
transform -1 0 7544 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _306_
timestamp 1704896540
transform 1 0 5520 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _307_
timestamp 1704896540
transform 1 0 6716 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _308_
timestamp 1704896540
transform -1 0 3772 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _309_
timestamp 1704896540
transform -1 0 7084 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _310_
timestamp 1704896540
transform 1 0 6072 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _311_
timestamp 1704896540
transform 1 0 8924 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _312_
timestamp 1704896540
transform 1 0 9384 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _313_
timestamp 1704896540
transform 1 0 10672 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _314_
timestamp 1704896540
transform -1 0 10396 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _315_
timestamp 1704896540
transform -1 0 11132 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _316_
timestamp 1704896540
transform 1 0 10488 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _317_
timestamp 1704896540
transform -1 0 14996 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _318_
timestamp 1704896540
transform 1 0 12696 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _319_
timestamp 1704896540
transform 1 0 14260 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _320_
timestamp 1704896540
transform 1 0 14720 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _321_
timestamp 1704896540
transform 1 0 13248 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _322_
timestamp 1704896540
transform -1 0 15180 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _323_
timestamp 1704896540
transform 1 0 11868 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _324_
timestamp 1704896540
transform 1 0 12512 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _325_
timestamp 1704896540
transform 1 0 13340 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _326_
timestamp 1704896540
transform 1 0 15548 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _327_
timestamp 1704896540
transform 1 0 13064 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _328_
timestamp 1704896540
transform 1 0 14076 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _329_
timestamp 1704896540
transform 1 0 12788 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _330_
timestamp 1704896540
transform 1 0 12696 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _331_
timestamp 1704896540
transform 1 0 13892 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _332_
timestamp 1704896540
transform 1 0 13800 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _333_
timestamp 1704896540
transform 1 0 13064 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _334_
timestamp 1704896540
transform -1 0 14996 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__mux4_1  _335_
timestamp 1704896540
transform 1 0 9200 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _336_
timestamp 1704896540
transform 1 0 10672 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _337_
timestamp 1704896540
transform 1 0 11500 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _338_
timestamp 1704896540
transform 1 0 12788 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _339_
timestamp 1704896540
transform 1 0 10672 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _340_
timestamp 1704896540
transform -1 0 11776 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4b_1  _341_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10120 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _342_
timestamp 1704896540
transform 1 0 10672 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _343_
timestamp 1704896540
transform 1 0 3772 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _344_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3404 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _345_
timestamp 1704896540
transform 1 0 2300 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _346_
timestamp 1704896540
transform 1 0 1564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _347_
timestamp 1704896540
transform 1 0 4508 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _348_
timestamp 1704896540
transform -1 0 3680 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _349_
timestamp 1704896540
transform 1 0 7452 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _350_
timestamp 1704896540
transform 1 0 7176 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _351_
timestamp 1704896540
transform 1 0 11592 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _352_
timestamp 1704896540
transform -1 0 11408 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _353_
timestamp 1704896540
transform -1 0 11408 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _354_
timestamp 1704896540
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _355_
timestamp 1704896540
transform 1 0 11684 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _356_
timestamp 1704896540
transform 1 0 11500 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _357_
timestamp 1704896540
transform 1 0 8372 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _358_
timestamp 1704896540
transform 1 0 8096 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _359_
timestamp 1704896540
transform 1 0 9844 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _360_
timestamp 1704896540
transform 1 0 11500 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _361_
timestamp 1704896540
transform 1 0 4692 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _362_
timestamp 1704896540
transform 1 0 4876 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _363_
timestamp 1704896540
transform 1 0 3864 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _364_
timestamp 1704896540
transform 1 0 3956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _365_
timestamp 1704896540
transform 1 0 6348 0 -1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _366_
timestamp 1704896540
transform 1 0 5612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _367_
timestamp 1704896540
transform 1 0 8004 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _368_
timestamp 1704896540
transform -1 0 7728 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _369_
timestamp 1704896540
transform -1 0 14996 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _370_
timestamp 1704896540
transform 1 0 15456 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _371_
timestamp 1704896540
transform 1 0 12144 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _372_
timestamp 1704896540
transform -1 0 11408 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _373_
timestamp 1704896540
transform 1 0 14076 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _374_
timestamp 1704896540
transform -1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _375_
timestamp 1704896540
transform 1 0 9476 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _376_
timestamp 1704896540
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_4  _377_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 8924 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _378_
timestamp 1704896540
transform 1 0 6256 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _379_
timestamp 1704896540
transform -1 0 6256 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _380_
timestamp 1704896540
transform -1 0 7728 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _381_
timestamp 1704896540
transform -1 0 7820 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _382_
timestamp 1704896540
transform -1 0 7728 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _383_
timestamp 1704896540
transform 1 0 7636 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _384_
timestamp 1704896540
transform -1 0 10212 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _385_
timestamp 1704896540
transform 1 0 10212 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _386_
timestamp 1704896540
transform -1 0 16284 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _387_
timestamp 1704896540
transform 1 0 16284 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _388_
timestamp 1704896540
transform 1 0 15456 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _389_
timestamp 1704896540
transform -1 0 15548 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _390_
timestamp 1704896540
transform 1 0 14812 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _391_
timestamp 1704896540
transform -1 0 14812 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _392_
timestamp 1704896540
transform 1 0 10580 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _393_
timestamp 1704896540
transform -1 0 9936 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and4b_1  _394_
timestamp 1704896540
transform 1 0 9844 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _395_
timestamp 1704896540
transform 1 0 10672 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _396_
timestamp 1704896540
transform 1 0 2116 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _397_
timestamp 1704896540
transform 1 0 1748 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _398_
timestamp 1704896540
transform 1 0 2208 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _399_
timestamp 1704896540
transform 1 0 1748 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _400_
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _401_
timestamp 1704896540
transform 1 0 2944 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _402_
timestamp 1704896540
transform -1 0 9384 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _403_
timestamp 1704896540
transform 1 0 9108 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _404_
timestamp 1704896540
transform -1 0 17388 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _405_
timestamp 1704896540
transform -1 0 17756 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _406_
timestamp 1704896540
transform 1 0 16652 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _407_
timestamp 1704896540
transform -1 0 16100 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _408_
timestamp 1704896540
transform -1 0 16560 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _409_
timestamp 1704896540
transform 1 0 16652 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _410_
timestamp 1704896540
transform 1 0 14996 0 1 4352
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _411_
timestamp 1704896540
transform 1 0 15180 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_4  _412_
timestamp 1704896540
transform -1 0 9660 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _413_
timestamp 1704896540
transform 1 0 2300 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _414_
timestamp 1704896540
transform 1 0 1932 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _415_
timestamp 1704896540
transform 1 0 2024 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _416_
timestamp 1704896540
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _417_
timestamp 1704896540
transform 1 0 2852 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _418_
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _419_
timestamp 1704896540
transform 1 0 7452 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _420_
timestamp 1704896540
transform 1 0 7268 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _421_
timestamp 1704896540
transform -1 0 16376 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _422_
timestamp 1704896540
transform 1 0 17572 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _423_
timestamp 1704896540
transform 1 0 16652 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _424_
timestamp 1704896540
transform -1 0 15824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _425_
timestamp 1704896540
transform -1 0 17296 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _426_
timestamp 1704896540
transform -1 0 17572 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _427_
timestamp 1704896540
transform -1 0 16468 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _428_
timestamp 1704896540
transform -1 0 16744 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or4b_1  _429_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 8832 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _430_
timestamp 1704896540
transform 1 0 8004 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _431_
timestamp 1704896540
transform 1 0 7084 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _432_
timestamp 1704896540
transform -1 0 6900 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _433_
timestamp 1704896540
transform 1 0 7268 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _434_
timestamp 1704896540
transform 1 0 7268 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _435_
timestamp 1704896540
transform -1 0 8280 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _436_
timestamp 1704896540
transform -1 0 8280 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _437_
timestamp 1704896540
transform 1 0 9936 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _438_
timestamp 1704896540
transform -1 0 9752 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _439_
timestamp 1704896540
transform -1 0 16376 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _440_
timestamp 1704896540
transform 1 0 17388 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _441_
timestamp 1704896540
transform -1 0 14904 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _442_
timestamp 1704896540
transform 1 0 14536 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _443_
timestamp 1704896540
transform 1 0 15180 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _444_
timestamp 1704896540
transform -1 0 14996 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _445_
timestamp 1704896540
transform -1 0 16192 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _446_
timestamp 1704896540
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and4bb_4  _447_
timestamp 1704896540
transform 1 0 8556 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _448_
timestamp 1704896540
transform 1 0 4232 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _449_
timestamp 1704896540
transform 1 0 3956 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _450_
timestamp 1704896540
transform 1 0 4232 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _451_
timestamp 1704896540
transform 1 0 3956 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _452_
timestamp 1704896540
transform -1 0 5520 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _453_
timestamp 1704896540
transform 1 0 5244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _454_
timestamp 1704896540
transform 1 0 8740 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _455_
timestamp 1704896540
transform 1 0 8464 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _456_
timestamp 1704896540
transform -1 0 12696 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _457_
timestamp 1704896540
transform 1 0 12420 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _458_
timestamp 1704896540
transform 1 0 11684 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _459_
timestamp 1704896540
transform 1 0 11500 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _460_
timestamp 1704896540
transform 1 0 11960 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _461_
timestamp 1704896540
transform 1 0 12052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _462_
timestamp 1704896540
transform 1 0 9108 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _463_
timestamp 1704896540
transform -1 0 9200 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _464_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 10856 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _465_
timestamp 1704896540
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _466_
timestamp 1704896540
transform 1 0 3772 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _467_
timestamp 1704896540
transform 1 0 2944 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _468_
timestamp 1704896540
transform 1 0 2944 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _469_
timestamp 1704896540
transform -1 0 2116 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _470_
timestamp 1704896540
transform 1 0 4508 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _471_
timestamp 1704896540
transform 1 0 4232 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _472_
timestamp 1704896540
transform 1 0 7176 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _473_
timestamp 1704896540
transform 1 0 6900 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _474_
timestamp 1704896540
transform -1 0 13984 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _475_
timestamp 1704896540
transform 1 0 13616 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _476_
timestamp 1704896540
transform 1 0 10948 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _477_
timestamp 1704896540
transform 1 0 10672 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _478_
timestamp 1704896540
transform -1 0 13064 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _479_
timestamp 1704896540
transform 1 0 12512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _480_
timestamp 1704896540
transform -1 0 8832 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _481_
timestamp 1704896540
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  _482_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3128 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _483_
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _484_
timestamp 1704896540
transform 1 0 4048 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _485_
timestamp 1704896540
transform 1 0 6900 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _486_
timestamp 1704896540
transform 1 0 11500 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _487_
timestamp 1704896540
transform 1 0 10304 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _488_
timestamp 1704896540
transform 1 0 11224 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _489_
timestamp 1704896540
transform 1 0 7360 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _490_
timestamp 1704896540
transform 1 0 4232 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _491_
timestamp 1704896540
transform 1 0 3496 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _492_
timestamp 1704896540
transform 1 0 5336 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _493_
timestamp 1704896540
transform 1 0 7912 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _494_
timestamp 1704896540
transform -1 0 15732 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _495_
timestamp 1704896540
transform 1 0 11684 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _496_
timestamp 1704896540
transform -1 0 14628 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _497_
timestamp 1704896540
transform 1 0 9016 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _498_
timestamp 1704896540
transform -1 0 7820 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _499_
timestamp 1704896540
transform -1 0 8096 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _500_
timestamp 1704896540
transform -1 0 7820 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _501_
timestamp 1704896540
transform 1 0 9108 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _502_
timestamp 1704896540
transform 1 0 16008 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _503_
timestamp 1704896540
transform 1 0 15548 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _504_
timestamp 1704896540
transform 1 0 14628 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _505_
timestamp 1704896540
transform -1 0 11408 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _506_
timestamp 1704896540
transform 1 0 1380 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _507_
timestamp 1704896540
transform 1 0 1380 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _508_
timestamp 1704896540
transform 1 0 2576 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _509_
timestamp 1704896540
transform 1 0 8924 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _510_
timestamp 1704896540
transform -1 0 17848 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _511_
timestamp 1704896540
transform -1 0 16560 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _512_
timestamp 1704896540
transform 1 0 16376 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _513_
timestamp 1704896540
transform 1 0 14720 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _514_
timestamp 1704896540
transform 1 0 1472 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _515_
timestamp 1704896540
transform 1 0 1564 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _516_
timestamp 1704896540
transform 1 0 2024 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _517_
timestamp 1704896540
transform 1 0 6900 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _518_
timestamp 1704896540
transform -1 0 17848 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _519_
timestamp 1704896540
transform -1 0 17848 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _520_
timestamp 1704896540
transform -1 0 17848 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _521_
timestamp 1704896540
transform -1 0 17388 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _522_
timestamp 1704896540
transform 1 0 6900 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _523_
timestamp 1704896540
transform 1 0 6532 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _524_
timestamp 1704896540
transform -1 0 8832 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _525_
timestamp 1704896540
transform 1 0 9752 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _526_
timestamp 1704896540
transform -1 0 16560 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _527_
timestamp 1704896540
transform -1 0 14904 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _528_
timestamp 1704896540
transform 1 0 14996 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _529_
timestamp 1704896540
transform -1 0 16560 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _530_
timestamp 1704896540
transform 1 0 3772 0 -1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _531_
timestamp 1704896540
transform 1 0 3588 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _532_
timestamp 1704896540
transform 1 0 4140 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _533_
timestamp 1704896540
transform 1 0 8004 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _534_
timestamp 1704896540
transform 1 0 11316 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _535_
timestamp 1704896540
transform 1 0 11224 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _536_
timestamp 1704896540
transform 1 0 11684 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _537_
timestamp 1704896540
transform 1 0 9200 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _538_
timestamp 1704896540
transform 1 0 2576 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _539_
timestamp 1704896540
transform 1 0 2116 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _540_
timestamp 1704896540
transform 1 0 4140 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _541_
timestamp 1704896540
transform 1 0 6440 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _542_
timestamp 1704896540
transform 1 0 13248 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _543_
timestamp 1704896540
transform 1 0 9936 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _544_
timestamp 1704896540
transform 1 0 11684 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _545_
timestamp 1704896540
transform 1 0 7820 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9476 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_0__f_clk
timestamp 1704896540
transform -1 0 6256 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_1__f_clk
timestamp 1704896540
transform 1 0 7360 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_2__f_clk
timestamp 1704896540
transform -1 0 6072 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_3__f_clk
timestamp 1704896540
transform -1 0 8832 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_4__f_clk
timestamp 1704896540
transform -1 0 13984 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_5__f_clk
timestamp 1704896540
transform 1 0 14352 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_6__f_clk
timestamp 1704896540
transform -1 0 13708 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_3_7__f_clk
timestamp 1704896540
transform 1 0 14720 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  clkload0
timestamp 1704896540
transform 1 0 4692 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkinvlp_2  clkload1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7636 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  clkload2
timestamp 1704896540
transform 1 0 4232 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__bufinv_16  clkload3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 12420 0 -1 6528
box -38 -48 2246 592
use sky130_fd_sc_hd__clkinvlp_2  clkload4
timestamp 1704896540
transform 1 0 14628 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  clkload5 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 11592 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  clkload6
timestamp 1704896540
transform 1 0 14444 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_3 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_15
timestamp 1704896540
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_35
timestamp 1704896540
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_47 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 5428 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_51
timestamp 1704896540
transform 1 0 5796 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1704896540
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_85
timestamp 1704896540
transform 1 0 8924 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_135
timestamp 1704896540
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1704896540
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_158 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 15640 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_166
timestamp 1704896540
transform 1 0 16376 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1704896540
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_181
timestamp 1704896540
transform 1 0 17756 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_52
timestamp 1704896540
transform 1 0 5888 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_113
timestamp 1704896540
transform 1 0 11500 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_163
timestamp 1704896540
transform 1 0 16100 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1704896540
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1704896540
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_181
timestamp 1704896540
transform 1 0 17756 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_29
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_33
timestamp 1704896540
transform 1 0 4140 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_62
timestamp 1704896540
transform 1 0 6808 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_72 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 7728 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_100
timestamp 1704896540
transform 1 0 10304 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_120
timestamp 1704896540
transform 1 0 12144 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_138
timestamp 1704896540
transform 1 0 13800 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_144
timestamp 1704896540
transform 1 0 14352 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_166
timestamp 1704896540
transform 1 0 16376 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1704896540
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1704896540
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_39
timestamp 1704896540
transform 1 0 4692 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_53
timestamp 1704896540
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_74
timestamp 1704896540
transform 1 0 7912 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_84
timestamp 1704896540
transform 1 0 8832 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_96
timestamp 1704896540
transform 1 0 9936 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_110
timestamp 1704896540
transform 1 0 11224 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_113
timestamp 1704896540
transform 1 0 11500 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_148
timestamp 1704896540
transform 1 0 14720 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_152
timestamp 1704896540
transform 1 0 15088 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_159
timestamp 1704896540
transform 1 0 15732 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_169
timestamp 1704896540
transform 1 0 16652 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_180
timestamp 1704896540
transform 1 0 17664 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_19
timestamp 1704896540
transform 1 0 2852 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_23
timestamp 1704896540
transform 1 0 3220 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_46
timestamp 1704896540
transform 1 0 5336 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_70
timestamp 1704896540
transform 1 0 7544 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_79
timestamp 1704896540
transform 1 0 8372 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1704896540
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_85
timestamp 1704896540
transform 1 0 8924 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_109
timestamp 1704896540
transform 1 0 11132 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_141
timestamp 1704896540
transform 1 0 14076 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_160
timestamp 1704896540
transform 1 0 15824 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_177
timestamp 1704896540
transform 1 0 17388 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_15
timestamp 1704896540
transform 1 0 2484 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_78
timestamp 1704896540
transform 1 0 8280 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_109
timestamp 1704896540
transform 1 0 11132 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_116
timestamp 1704896540
transform 1 0 11776 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_124
timestamp 1704896540
transform 1 0 12512 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_164
timestamp 1704896540
transform 1 0 16192 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_181
timestamp 1704896540
transform 1 0 17756 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_15
timestamp 1704896540
transform 1 0 2484 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_23
timestamp 1704896540
transform 1 0 3220 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_46
timestamp 1704896540
transform 1 0 5336 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_66
timestamp 1704896540
transform 1 0 7176 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_93
timestamp 1704896540
transform 1 0 9660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_101
timestamp 1704896540
transform 1 0 10396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_116
timestamp 1704896540
transform 1 0 11776 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_120
timestamp 1704896540
transform 1 0 12144 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_136
timestamp 1704896540
transform 1 0 13616 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_156
timestamp 1704896540
transform 1 0 15456 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_170
timestamp 1704896540
transform 1 0 16744 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_18
timestamp 1704896540
transform 1 0 2760 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_38
timestamp 1704896540
transform 1 0 4600 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_78
timestamp 1704896540
transform 1 0 8280 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_84
timestamp 1704896540
transform 1 0 8832 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_88
timestamp 1704896540
transform 1 0 9200 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_100
timestamp 1704896540
transform 1 0 10304 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_113
timestamp 1704896540
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_147
timestamp 1704896540
transform 1 0 14628 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_3
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_9
timestamp 1704896540
transform 1 0 1932 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1704896540
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_49
timestamp 1704896540
transform 1 0 5612 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_85
timestamp 1704896540
transform 1 0 8924 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_118
timestamp 1704896540
transform 1 0 11960 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_154
timestamp 1704896540
transform 1 0 15272 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_164
timestamp 1704896540
transform 1 0 16192 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_57
timestamp 1704896540
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_121
timestamp 1704896540
transform 1 0 12236 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_151
timestamp 1704896540
transform 1 0 14996 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_169
timestamp 1704896540
transform 1 0 16652 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1704896540
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_37
timestamp 1704896540
transform 1 0 4508 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_48
timestamp 1704896540
transform 1 0 5520 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_60
timestamp 1704896540
transform 1 0 6624 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_78
timestamp 1704896540
transform 1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1704896540
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_97
timestamp 1704896540
transform 1 0 10028 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_103
timestamp 1704896540
transform 1 0 10580 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_110
timestamp 1704896540
transform 1 0 11224 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_118
timestamp 1704896540
transform 1 0 11960 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_125
timestamp 1704896540
transform 1 0 12604 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_141
timestamp 1704896540
transform 1 0 14076 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_164
timestamp 1704896540
transform 1 0 16192 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_19
timestamp 1704896540
transform 1 0 2852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_29
timestamp 1704896540
transform 1 0 3772 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_34
timestamp 1704896540
transform 1 0 4232 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_57
timestamp 1704896540
transform 1 0 6348 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_72
timestamp 1704896540
transform 1 0 7728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_94
timestamp 1704896540
transform 1 0 9752 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_103
timestamp 1704896540
transform 1 0 10580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_110
timestamp 1704896540
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_113
timestamp 1704896540
transform 1 0 11500 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_117
timestamp 1704896540
transform 1 0 11868 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_127
timestamp 1704896540
transform 1 0 12788 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_137
timestamp 1704896540
transform 1 0 13708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_147
timestamp 1704896540
transform 1 0 14628 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_162
timestamp 1704896540
transform 1 0 16008 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1704896540
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_3
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1704896540
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_113
timestamp 1704896540
transform 1 0 11500 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1704896540
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_147
timestamp 1704896540
transform 1 0 14628 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_179
timestamp 1704896540
transform 1 0 17572 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_3
timestamp 1704896540
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_22
timestamp 1704896540
transform 1 0 3128 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_50
timestamp 1704896540
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_63
timestamp 1704896540
transform 1 0 6900 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_78
timestamp 1704896540
transform 1 0 8280 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_93
timestamp 1704896540
transform 1 0 9660 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_103
timestamp 1704896540
transform 1 0 10580 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1704896540
transform 1 0 11224 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_122
timestamp 1704896540
transform 1 0 12328 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_150
timestamp 1704896540
transform 1 0 14904 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_158
timestamp 1704896540
transform 1 0 15640 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_177
timestamp 1704896540
transform 1 0 17388 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_181
timestamp 1704896540
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_11
timestamp 1704896540
transform 1 0 2116 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_21
timestamp 1704896540
transform 1 0 3036 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1704896540
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 1704896540
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 1704896540
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 1704896540
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_65
timestamp 1704896540
transform 1 0 7084 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_73
timestamp 1704896540
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1704896540
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_85
timestamp 1704896540
transform 1 0 8924 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_93
timestamp 1704896540
transform 1 0 9660 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_131
timestamp 1704896540
transform 1 0 13156 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_158
timestamp 1704896540
transform 1 0 15640 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_163
timestamp 1704896540
transform 1 0 16100 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_179
timestamp 1704896540
transform 1 0 17572 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_19
timestamp 1704896540
transform 1 0 2852 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_23
timestamp 1704896540
transform 1 0 3220 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_41
timestamp 1704896540
transform 1 0 4876 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_57
timestamp 1704896540
transform 1 0 6348 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1704896540
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_113
timestamp 1704896540
transform 1 0 11500 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_149
timestamp 1704896540
transform 1 0 14812 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_29
timestamp 1704896540
transform 1 0 3772 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_57
timestamp 1704896540
transform 1 0 6348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_66
timestamp 1704896540
transform 1 0 7176 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_85
timestamp 1704896540
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_134
timestamp 1704896540
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_141
timestamp 1704896540
transform 1 0 14076 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_147
timestamp 1704896540
transform 1 0 14628 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 1704896540
transform 1 0 1380 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_21
timestamp 1704896540
transform 1 0 3036 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 1704896540
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1704896540
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_65
timestamp 1704896540
transform 1 0 7084 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_77
timestamp 1704896540
transform 1 0 8188 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_100
timestamp 1704896540
transform 1 0 10304 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_116
timestamp 1704896540
transform 1 0 11776 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_124
timestamp 1704896540
transform 1 0 12512 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_131
timestamp 1704896540
transform 1 0 13156 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_149
timestamp 1704896540
transform 1 0 14812 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_181
timestamp 1704896540
transform 1 0 17756 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_12
timestamp 1704896540
transform 1 0 2208 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_26
timestamp 1704896540
transform 1 0 3496 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_29
timestamp 1704896540
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_74
timestamp 1704896540
transform 1 0 7912 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_78
timestamp 1704896540
transform 1 0 8280 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_82
timestamp 1704896540
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_88
timestamp 1704896540
transform 1 0 9200 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_96
timestamp 1704896540
transform 1 0 9936 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_112
timestamp 1704896540
transform 1 0 11408 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_124
timestamp 1704896540
transform 1 0 12512 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 1704896540
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 1704896540
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_141
timestamp 1704896540
transform 1 0 14076 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_151
timestamp 1704896540
transform 1 0 14996 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_9
timestamp 1704896540
transform 1 0 1932 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_45
timestamp 1704896540
transform 1 0 5244 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_57
timestamp 1704896540
transform 1 0 6348 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_87
timestamp 1704896540
transform 1 0 9108 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_102
timestamp 1704896540
transform 1 0 10488 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_113
timestamp 1704896540
transform 1 0 11500 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_148
timestamp 1704896540
transform 1 0 14720 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_180
timestamp 1704896540
transform 1 0 17664 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_29
timestamp 1704896540
transform 1 0 3772 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_33
timestamp 1704896540
transform 1 0 4140 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_54
timestamp 1704896540
transform 1 0 6072 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 1704896540
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 1704896540
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 1704896540
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_85
timestamp 1704896540
transform 1 0 8924 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_91
timestamp 1704896540
transform 1 0 9476 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_109
timestamp 1704896540
transform 1 0 11132 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_135
timestamp 1704896540
transform 1 0 13524 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1704896540
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_141
timestamp 1704896540
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_177
timestamp 1704896540
transform 1 0 17388 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_3
timestamp 1704896540
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_10
timestamp 1704896540
transform 1 0 2024 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_16
timestamp 1704896540
transform 1 0 2576 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_25
timestamp 1704896540
transform 1 0 3404 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_33
timestamp 1704896540
transform 1 0 4140 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_40
timestamp 1704896540
transform 1 0 4784 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_44
timestamp 1704896540
transform 1 0 5152 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 1704896540
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 1704896540
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_65
timestamp 1704896540
transform 1 0 7084 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_78
timestamp 1704896540
transform 1 0 8280 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_90
timestamp 1704896540
transform 1 0 9384 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_102
timestamp 1704896540
transform 1 0 10488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_110
timestamp 1704896540
transform 1 0 11224 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_113
timestamp 1704896540
transform 1 0 11500 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_126
timestamp 1704896540
transform 1 0 12696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_130
timestamp 1704896540
transform 1 0 13064 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_137
timestamp 1704896540
transform 1 0 13708 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_141
timestamp 1704896540
transform 1 0 14076 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_166
timestamp 1704896540
transform 1 0 16376 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_169
timestamp 1704896540
transform 1 0 16652 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_7
timestamp 1704896540
transform 1 0 1748 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_12
timestamp 1704896540
transform 1 0 2208 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_22
timestamp 1704896540
transform 1 0 3128 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 1704896540
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 1704896540
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_53
timestamp 1704896540
transform 1 0 5980 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_60
timestamp 1704896540
transform 1 0 6624 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_109
timestamp 1704896540
transform 1 0 11132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_113
timestamp 1704896540
transform 1 0 11500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_137
timestamp 1704896540
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_153
timestamp 1704896540
transform 1 0 15180 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_3
timestamp 1704896540
transform 1 0 1380 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_28
timestamp 1704896540
transform 1 0 3680 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_34
timestamp 1704896540
transform 1 0 4232 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_90
timestamp 1704896540
transform 1 0 9384 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_108
timestamp 1704896540
transform 1 0 11040 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_129
timestamp 1704896540
transform 1 0 12972 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_151
timestamp 1704896540
transform 1 0 14996 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_155
timestamp 1704896540
transform 1 0 15364 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_169
timestamp 1704896540
transform 1 0 16652 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_7
timestamp 1704896540
transform 1 0 1748 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_19
timestamp 1704896540
transform 1 0 2852 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_38
timestamp 1704896540
transform 1 0 4600 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_61
timestamp 1704896540
transform 1 0 6716 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_70
timestamp 1704896540
transform 1 0 7544 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_82
timestamp 1704896540
transform 1 0 8648 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_106
timestamp 1704896540
transform 1 0 10856 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_118
timestamp 1704896540
transform 1 0 11960 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_132
timestamp 1704896540
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 1704896540
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_15
timestamp 1704896540
transform 1 0 2484 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_21
timestamp 1704896540
transform 1 0 3036 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_46
timestamp 1704896540
transform 1 0 5336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_54
timestamp 1704896540
transform 1 0 6072 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_57
timestamp 1704896540
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_65
timestamp 1704896540
transform 1 0 7084 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_78
timestamp 1704896540
transform 1 0 8280 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_102
timestamp 1704896540
transform 1 0 10488 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_116
timestamp 1704896540
transform 1 0 11776 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_138
timestamp 1704896540
transform 1 0 13800 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_150
timestamp 1704896540
transform 1 0 14904 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_165
timestamp 1704896540
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_177
timestamp 1704896540
transform 1 0 17388 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_7
timestamp 1704896540
transform 1 0 1748 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_19
timestamp 1704896540
transform 1 0 2852 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_23
timestamp 1704896540
transform 1 0 3220 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1704896540
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_38
timestamp 1704896540
transform 1 0 4600 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_56
timestamp 1704896540
transform 1 0 6256 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_62
timestamp 1704896540
transform 1 0 6808 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_79
timestamp 1704896540
transform 1 0 8372 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 1704896540
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_93
timestamp 1704896540
transform 1 0 9660 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_99
timestamp 1704896540
transform 1 0 10212 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_116
timestamp 1704896540
transform 1 0 11776 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_138
timestamp 1704896540
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 1704896540
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_153
timestamp 1704896540
transform 1 0 15180 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_181
timestamp 1704896540
transform 1 0 17756 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1704896540
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_15
timestamp 1704896540
transform 1 0 2484 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_32
timestamp 1704896540
transform 1 0 4048 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_50
timestamp 1704896540
transform 1 0 5704 0 -1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_73
timestamp 1704896540
transform 1 0 7820 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_85
timestamp 1704896540
transform 1 0 8924 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_89
timestamp 1704896540
transform 1 0 9292 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_102
timestamp 1704896540
transform 1 0 10488 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 1704896540
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 1704896540
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_137
timestamp 1704896540
transform 1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_141
timestamp 1704896540
transform 1 0 14076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_151
timestamp 1704896540
transform 1 0 14996 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_163
timestamp 1704896540
transform 1 0 16100 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1704896540
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 1704896540
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_181
timestamp 1704896540
transform 1 0 17756 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 1704896540
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 1704896540
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 1704896540
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_29
timestamp 1704896540
transform 1 0 3772 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_44
timestamp 1704896540
transform 1 0 5152 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_65
timestamp 1704896540
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_85
timestamp 1704896540
transform 1 0 8924 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_103
timestamp 1704896540
transform 1 0 10580 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_116
timestamp 1704896540
transform 1 0 11776 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_129
timestamp 1704896540
transform 1 0 12972 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_141
timestamp 1704896540
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_167
timestamp 1704896540
transform 1 0 16468 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_179
timestamp 1704896540
transform 1 0 17572 0 1 17408
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 1704896540
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 1704896540
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 1704896540
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 1704896540
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 1704896540
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 1704896540
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_57
timestamp 1704896540
transform 1 0 6348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_113
timestamp 1704896540
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_131
timestamp 1704896540
transform 1 0 13156 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_159
timestamp 1704896540
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1704896540
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 1704896540
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_181
timestamp 1704896540
transform 1 0 17756 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 1704896540
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 1704896540
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 1704896540
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 1704896540
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1704896540
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_53
timestamp 1704896540
transform 1 0 5980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_57
timestamp 1704896540
transform 1 0 6348 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_66
timestamp 1704896540
transform 1 0 7176 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_107
timestamp 1704896540
transform 1 0 10948 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_121
timestamp 1704896540
transform 1 0 12236 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1704896540
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 1704896540
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 1704896540
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_165
timestamp 1704896540
transform 1 0 16284 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_169
timestamp 1704896540
transform 1 0 16652 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_181
timestamp 1704896540
transform 1 0 17756 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5704 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1704896540
transform -1 0 5336 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1704896540
transform -1 0 9660 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1704896540
transform -1 0 13800 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1704896540
transform -1 0 17388 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1704896540
transform -1 0 5796 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1704896540
transform -1 0 3680 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1704896540
transform -1 0 11408 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1704896540
transform -1 0 3496 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1704896540
transform -1 0 9660 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1704896540
transform -1 0 13616 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1704896540
transform -1 0 7912 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1704896540
transform -1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1704896540
transform -1 0 13432 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 1704896540
transform -1 0 12236 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 1704896540
transform -1 0 6256 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 1704896540
transform -1 0 12144 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 1704896540
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 1704896540
transform -1 0 4508 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 1704896540
transform -1 0 8832 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 1704896540
transform -1 0 17572 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 1704896540
transform -1 0 5796 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 1704896540
transform -1 0 13432 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 1704896540
transform -1 0 10304 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 1704896540
transform -1 0 5980 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 1704896540
transform -1 0 4876 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold27
timestamp 1704896540
transform -1 0 11408 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold28
timestamp 1704896540
transform -1 0 9660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold29
timestamp 1704896540
transform -1 0 13524 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold30
timestamp 1704896540
transform 1 0 6992 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold31
timestamp 1704896540
transform -1 0 6256 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold32
timestamp 1704896540
transform -1 0 13892 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold33
timestamp 1704896540
transform 1 0 6900 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold34
timestamp 1704896540
transform -1 0 10948 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold35
timestamp 1704896540
transform -1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold36
timestamp 1704896540
transform -1 0 3404 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold37
timestamp 1704896540
transform -1 0 16468 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold38
timestamp 1704896540
transform -1 0 16376 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold39
timestamp 1704896540
transform 1 0 1564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold40
timestamp 1704896540
transform -1 0 15640 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold41
timestamp 1704896540
transform 1 0 10488 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold42
timestamp 1704896540
transform 1 0 15824 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold43
timestamp 1704896540
transform -1 0 9108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold44
timestamp 1704896540
transform -1 0 8464 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold45
timestamp 1704896540
transform -1 0 4876 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold46
timestamp 1704896540
transform -1 0 17756 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold47
timestamp 1704896540
transform -1 0 15456 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold48
timestamp 1704896540
transform -1 0 5336 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold49
timestamp 1704896540
transform 1 0 16836 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold50
timestamp 1704896540
transform 1 0 5520 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold51
timestamp 1704896540
transform -1 0 11132 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold52
timestamp 1704896540
transform -1 0 17664 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold53
timestamp 1704896540
transform -1 0 16560 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold54
timestamp 1704896540
transform -1 0 17848 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold55
timestamp 1704896540
transform -1 0 6256 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold56
timestamp 1704896540
transform -1 0 17388 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold57
timestamp 1704896540
transform -1 0 15640 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold58
timestamp 1704896540
transform -1 0 9108 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold59
timestamp 1704896540
transform -1 0 17388 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold60
timestamp 1704896540
transform -1 0 8832 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold61
timestamp 1704896540
transform 1 0 6624 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold62
timestamp 1704896540
transform -1 0 17388 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold63
timestamp 1704896540
transform -1 0 11500 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold64
timestamp 1704896540
transform 1 0 14996 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 17848 0 1 5440
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 1704896540
transform -1 0 17848 0 -1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input3
timestamp 1704896540
transform 1 0 1380 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1704896540
transform -1 0 17848 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input5
timestamp 1704896540
transform 1 0 16928 0 -1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1704896540
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input7 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 9292 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 1704896540
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1704896540
transform 1 0 1380 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1704896540
transform 1 0 3956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1704896540
transform -1 0 8832 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input12
timestamp 1704896540
transform -1 0 17848 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input13
timestamp 1704896540
transform -1 0 17848 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1704896540
transform -1 0 17848 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input15
timestamp 1704896540
transform 1 0 13156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1704896540
transform 1 0 11500 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1704896540
transform 1 0 10488 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input18
timestamp 1704896540
transform -1 0 8832 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  output19
timestamp 1704896540
transform -1 0 1748 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output20
timestamp 1704896540
transform -1 0 2116 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output21
timestamp 1704896540
transform 1 0 5888 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1704896540
transform -1 0 9936 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output23
timestamp 1704896540
transform 1 0 17480 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1704896540
transform -1 0 12880 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1704896540
transform 1 0 17480 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output26
timestamp 1704896540
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output27
timestamp 1704896540
transform -1 0 1748 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1704896540
transform -1 0 1748 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output29
timestamp 1704896540
transform 1 0 6532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1704896540
transform 1 0 9660 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output31
timestamp 1704896540
transform 1 0 17480 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output32
timestamp 1704896540
transform 1 0 16744 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output33
timestamp 1704896540
transform 1 0 17388 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output34
timestamp 1704896540
transform 1 0 12420 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_31
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 18124 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_32
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_33
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_34
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 18124 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_35
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 18124 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_36
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 18124 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_37
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 18124 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_38
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 18124 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_39
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 18124 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_40
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_41
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_42
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 18124 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_43
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 18124 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Left_44
timestamp 1704896540
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_13_Right_13
timestamp 1704896540
transform -1 0 18124 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Left_45
timestamp 1704896540
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_14_Right_14
timestamp 1704896540
transform -1 0 18124 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Left_46
timestamp 1704896540
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_15_Right_15
timestamp 1704896540
transform -1 0 18124 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Left_47
timestamp 1704896540
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_16_Right_16
timestamp 1704896540
transform -1 0 18124 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Left_48
timestamp 1704896540
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_17_Right_17
timestamp 1704896540
transform -1 0 18124 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Left_49
timestamp 1704896540
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_18_Right_18
timestamp 1704896540
transform -1 0 18124 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Left_50
timestamp 1704896540
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_19_Right_19
timestamp 1704896540
transform -1 0 18124 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Left_51
timestamp 1704896540
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_20_Right_20
timestamp 1704896540
transform -1 0 18124 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Left_52
timestamp 1704896540
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_21_Right_21
timestamp 1704896540
transform -1 0 18124 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Left_53
timestamp 1704896540
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_22_Right_22
timestamp 1704896540
transform -1 0 18124 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Left_54
timestamp 1704896540
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_23_Right_23
timestamp 1704896540
transform -1 0 18124 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Left_55
timestamp 1704896540
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_24_Right_24
timestamp 1704896540
transform -1 0 18124 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Left_56
timestamp 1704896540
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_25_Right_25
timestamp 1704896540
transform -1 0 18124 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Left_57
timestamp 1704896540
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_26_Right_26
timestamp 1704896540
transform -1 0 18124 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Left_58
timestamp 1704896540
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_27_Right_27
timestamp 1704896540
transform -1 0 18124 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Left_59
timestamp 1704896540
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_28_Right_28
timestamp 1704896540
transform -1 0 18124 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Left_60
timestamp 1704896540
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_29_Right_29
timestamp 1704896540
transform -1 0 18124 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Left_61
timestamp 1704896540
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_30_Right_30
timestamp 1704896540
transform -1 0 18124 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_62 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_63
timestamp 1704896540
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_64
timestamp 1704896540
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_65
timestamp 1704896540
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_66
timestamp 1704896540
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_67
timestamp 1704896540
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_68
timestamp 1704896540
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_69
timestamp 1704896540
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_1_70
timestamp 1704896540
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_71
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_72
timestamp 1704896540
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_73
timestamp 1704896540
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_74
timestamp 1704896540
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_75
timestamp 1704896540
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_3_76
timestamp 1704896540
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_77
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_78
timestamp 1704896540
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_79
timestamp 1704896540
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_80
timestamp 1704896540
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_81
timestamp 1704896540
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_5_82
timestamp 1704896540
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_83
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_84
timestamp 1704896540
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_85
timestamp 1704896540
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_86
timestamp 1704896540
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_87
timestamp 1704896540
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_7_88
timestamp 1704896540
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_89
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_90
timestamp 1704896540
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_91
timestamp 1704896540
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_92
timestamp 1704896540
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_93
timestamp 1704896540
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_9_94
timestamp 1704896540
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_95
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_96
timestamp 1704896540
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_97
timestamp 1704896540
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_98
timestamp 1704896540
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_99
timestamp 1704896540
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_11_100
timestamp 1704896540
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_101
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_102
timestamp 1704896540
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_103
timestamp 1704896540
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_104
timestamp 1704896540
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_105
timestamp 1704896540
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_13_106
timestamp 1704896540
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_107
timestamp 1704896540
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_108
timestamp 1704896540
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_14_109
timestamp 1704896540
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_110
timestamp 1704896540
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_111
timestamp 1704896540
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_15_112
timestamp 1704896540
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_113
timestamp 1704896540
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_114
timestamp 1704896540
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_16_115
timestamp 1704896540
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_116
timestamp 1704896540
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_117
timestamp 1704896540
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_17_118
timestamp 1704896540
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_119
timestamp 1704896540
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_120
timestamp 1704896540
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_18_121
timestamp 1704896540
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_122
timestamp 1704896540
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_123
timestamp 1704896540
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_19_124
timestamp 1704896540
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_125
timestamp 1704896540
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_126
timestamp 1704896540
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_20_127
timestamp 1704896540
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_128
timestamp 1704896540
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_129
timestamp 1704896540
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_21_130
timestamp 1704896540
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_131
timestamp 1704896540
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_132
timestamp 1704896540
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_22_133
timestamp 1704896540
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_134
timestamp 1704896540
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_135
timestamp 1704896540
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_23_136
timestamp 1704896540
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_137
timestamp 1704896540
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_138
timestamp 1704896540
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_24_139
timestamp 1704896540
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_140
timestamp 1704896540
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_141
timestamp 1704896540
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_25_142
timestamp 1704896540
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_143
timestamp 1704896540
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_144
timestamp 1704896540
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_26_145
timestamp 1704896540
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_146
timestamp 1704896540
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_147
timestamp 1704896540
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_27_148
timestamp 1704896540
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_149
timestamp 1704896540
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_150
timestamp 1704896540
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_28_151
timestamp 1704896540
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_152
timestamp 1704896540
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_153
timestamp 1704896540
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_29_154
timestamp 1704896540
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_155
timestamp 1704896540
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_156
timestamp 1704896540
transform 1 0 6256 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_157
timestamp 1704896540
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_158
timestamp 1704896540
transform 1 0 11408 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_159
timestamp 1704896540
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_30_160
timestamp 1704896540
transform 1 0 16560 0 1 18496
box -38 -48 130 592
<< labels >>
flabel metal4 s 3731 2128 4051 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 7986 2128 8306 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 12241 2128 12561 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 16496 2128 16816 19088 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 4784 18172 5104 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 9000 18172 9320 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 13216 18172 13536 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 17432 18172 17752 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 3071 2128 3391 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 7326 2128 7646 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 11581 2128 11901 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 15836 2128 16156 19088 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 4124 18172 4444 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 8340 18172 8660 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 12556 18172 12876 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 16772 18172 17092 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 17688 800 17808 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 0 14968 800 15088 0 FreeSans 480 0 0 0 readData1[0]
port 3 nsew signal output
flabel metal3 s 0 9528 800 9648 0 FreeSans 480 0 0 0 readData1[1]
port 4 nsew signal output
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 readData1[2]
port 5 nsew signal output
flabel metal2 s 9678 20613 9734 21413 0 FreeSans 224 90 0 0 readData1[3]
port 6 nsew signal output
flabel metal3 s 18469 15648 19269 15768 0 FreeSans 480 0 0 0 readData1[4]
port 7 nsew signal output
flabel metal2 s 12898 20613 12954 21413 0 FreeSans 224 90 0 0 readData1[5]
port 8 nsew signal output
flabel metal3 s 18469 5448 19269 5568 0 FreeSans 480 0 0 0 readData1[6]
port 9 nsew signal output
flabel metal2 s 11610 0 11666 800 0 FreeSans 224 90 0 0 readData1[7]
port 10 nsew signal output
flabel metal3 s 0 14288 800 14408 0 FreeSans 480 0 0 0 readData2[0]
port 11 nsew signal output
flabel metal3 s 0 10208 800 10328 0 FreeSans 480 0 0 0 readData2[1]
port 12 nsew signal output
flabel metal2 s 7102 0 7158 800 0 FreeSans 224 90 0 0 readData2[2]
port 13 nsew signal output
flabel metal2 s 10322 20613 10378 21413 0 FreeSans 224 90 0 0 readData2[3]
port 14 nsew signal output
flabel metal3 s 18469 14968 19269 15088 0 FreeSans 480 0 0 0 readData2[4]
port 15 nsew signal output
flabel metal3 s 18469 14288 19269 14408 0 FreeSans 480 0 0 0 readData2[5]
port 16 nsew signal output
flabel metal3 s 18469 4768 19269 4888 0 FreeSans 480 0 0 0 readData2[6]
port 17 nsew signal output
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 readData2[7]
port 18 nsew signal output
flabel metal3 s 18469 6128 19269 6248 0 FreeSans 480 0 0 0 readReg1[0]
port 19 nsew signal input
flabel metal3 s 18469 7488 19269 7608 0 FreeSans 480 0 0 0 readReg1[1]
port 20 nsew signal input
flabel metal3 s 0 12928 800 13048 0 FreeSans 480 0 0 0 readReg1[2]
port 21 nsew signal input
flabel metal3 s 18469 6808 19269 6928 0 FreeSans 480 0 0 0 readReg2[0]
port 22 nsew signal input
flabel metal3 s 18469 8168 19269 8288 0 FreeSans 480 0 0 0 readReg2[1]
port 23 nsew signal input
flabel metal3 s 0 12248 800 12368 0 FreeSans 480 0 0 0 readReg2[2]
port 24 nsew signal input
flabel metal2 s 9034 0 9090 800 0 FreeSans 224 90 0 0 regWrite
port 25 nsew signal input
flabel metal3 s 0 16328 800 16448 0 FreeSans 480 0 0 0 writeData[0]
port 26 nsew signal input
flabel metal3 s 0 10888 800 11008 0 FreeSans 480 0 0 0 writeData[1]
port 27 nsew signal input
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 writeData[2]
port 28 nsew signal input
flabel metal2 s 9034 20613 9090 21413 0 FreeSans 224 90 0 0 writeData[3]
port 29 nsew signal input
flabel metal3 s 18469 12928 19269 13048 0 FreeSans 480 0 0 0 writeData[4]
port 30 nsew signal input
flabel metal3 s 18469 10208 19269 10328 0 FreeSans 480 0 0 0 writeData[5]
port 31 nsew signal input
flabel metal3 s 18469 3408 19269 3528 0 FreeSans 480 0 0 0 writeData[6]
port 32 nsew signal input
flabel metal2 s 12254 0 12310 800 0 FreeSans 224 90 0 0 writeData[7]
port 33 nsew signal input
flabel metal2 s 9678 0 9734 800 0 FreeSans 224 90 0 0 writeReg[0]
port 34 nsew signal input
flabel metal2 s 10322 0 10378 800 0 FreeSans 224 90 0 0 writeReg[1]
port 35 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 writeReg[2]
port 36 nsew signal input
rlabel metal1 9614 18496 9614 18496 0 VGND
rlabel metal1 9614 19040 9614 19040 0 VPWR
rlabel metal2 3450 15878 3450 15878 0 _000_
rlabel via1 1697 8466 1697 8466 0 _001_
rlabel via1 4365 5270 4365 5270 0 _002_
rlabel metal2 7222 16354 7222 16354 0 _003_
rlabel metal1 11576 15062 11576 15062 0 _004_
rlabel metal2 11546 16354 11546 16354 0 _005_
rlabel metal1 11438 4522 11438 4522 0 _006_
rlabel metal1 7958 4794 7958 4794 0 _007_
rlabel metal1 4733 17238 4733 17238 0 _008_
rlabel metal1 3818 8602 3818 8602 0 _009_
rlabel metal2 5658 3298 5658 3298 0 _010_
rlabel metal1 8080 18326 8080 18326 0 _011_
rlabel via1 15414 17646 15414 17646 0 _012_
rlabel metal1 11904 18258 11904 18258 0 _013_
rlabel via1 14310 3026 14310 3026 0 _014_
rlabel via1 9333 2414 9333 2414 0 _015_
rlabel metal1 6858 17170 6858 17170 0 _016_
rlabel via1 7778 8942 7778 8942 0 _017_
rlabel metal1 7600 3026 7600 3026 0 _018_
rlabel metal2 10258 17442 10258 17442 0 _019_
rlabel metal2 16330 15266 16330 15266 0 _020_
rlabel metal1 15670 16490 15670 16490 0 _021_
rlabel metal1 14842 3094 14842 3094 0 _022_
rlabel metal1 10492 3094 10492 3094 0 _023_
rlabel via1 1697 13294 1697 13294 0 _024_
rlabel metal1 1743 10710 1743 10710 0 _025_
rlabel metal1 2944 4794 2944 4794 0 _026_
rlabel via1 9241 14382 9241 14382 0 _027_
rlabel metal2 17710 12002 17710 12002 0 _028_
rlabel metal1 16146 10234 16146 10234 0 _029_
rlabel metal1 16790 6426 16790 6426 0 _030_
rlabel metal1 15129 5270 15129 5270 0 _031_
rlabel metal1 1886 14586 1886 14586 0 _032_
rlabel via1 1881 11730 1881 11730 0 _033_
rlabel metal2 2530 6562 2530 6562 0 _034_
rlabel metal1 7263 15062 7263 15062 0 _035_
rlabel viali 17530 14382 17530 14382 0 _036_
rlabel metal1 16656 11050 16656 11050 0 _037_
rlabel via1 17530 7786 17530 7786 0 _038_
rlabel via1 17070 4522 17070 4522 0 _039_
rlabel metal1 7022 12886 7022 12886 0 _040_
rlabel metal1 7084 10234 7084 10234 0 _041_
rlabel metal2 8418 6562 8418 6562 0 _042_
rlabel metal1 9874 11050 9874 11050 0 _043_
rlabel metal1 16851 12886 16851 12886 0 _044_
rlabel via1 14586 9622 14586 9622 0 _045_
rlabel metal1 15118 8874 15118 8874 0 _046_
rlabel metal1 16340 7378 16340 7378 0 _047_
rlabel via1 4089 12818 4089 12818 0 _048_
rlabel metal1 3956 11322 3956 11322 0 _049_
rlabel metal1 4871 6766 4871 6766 0 _050_
rlabel metal1 8413 10710 8413 10710 0 _051_
rlabel metal2 12466 13498 12466 13498 0 _052_
rlabel metal1 11909 11118 11909 11118 0 _053_
rlabel metal1 12047 8874 12047 8874 0 _054_
rlabel metal2 9154 6902 9154 6902 0 _055_
rlabel metal1 2944 16762 2944 16762 0 _056_
rlabel metal1 2238 8874 2238 8874 0 _057_
rlabel metal1 4354 3094 4354 3094 0 _058_
rlabel via1 6757 18258 6757 18258 0 _059_
rlabel metal1 13611 18326 13611 18326 0 _060_
rlabel metal2 10718 18054 10718 18054 0 _061_
rlabel via1 12001 3026 12001 3026 0 _062_
rlabel metal1 8551 3094 8551 3094 0 _063_
rlabel metal1 13202 13940 13202 13940 0 _064_
rlabel metal2 12742 5338 12742 5338 0 _065_
rlabel metal1 6670 11220 6670 11220 0 _066_
rlabel via1 14196 12818 14196 12818 0 _067_
rlabel metal1 6716 14994 6716 14994 0 _068_
rlabel metal1 6670 13872 6670 13872 0 _069_
rlabel metal1 12742 11730 12742 11730 0 _070_
rlabel via1 6509 13906 6509 13906 0 _071_
rlabel metal1 15180 13158 15180 13158 0 _072_
rlabel metal1 4094 12614 4094 12614 0 _073_
rlabel metal1 6486 14042 6486 14042 0 _074_
rlabel metal2 6578 9248 6578 9248 0 _075_
rlabel metal1 5750 10506 5750 10506 0 _076_
rlabel metal1 6325 11118 6325 11118 0 _077_
rlabel metal1 4784 11050 4784 11050 0 _078_
rlabel metal1 6440 9554 6440 9554 0 _079_
rlabel metal1 7636 5338 7636 5338 0 _080_
rlabel metal1 6946 6154 6946 6154 0 _081_
rlabel metal1 6555 6766 6555 6766 0 _082_
rlabel metal2 4554 6562 4554 6562 0 _083_
rlabel metal2 6854 6154 6854 6154 0 _084_
rlabel metal2 10350 15436 10350 15436 0 _085_
rlabel metal1 10166 12784 10166 12784 0 _086_
rlabel metal1 10511 12818 10511 12818 0 _087_
rlabel metal1 9890 12886 9890 12886 0 _088_
rlabel metal2 10442 13787 10442 13787 0 _089_
rlabel metal2 14306 14620 14306 14620 0 _090_
rlabel metal1 13846 12342 13846 12342 0 _091_
rlabel via1 14492 12818 14492 12818 0 _092_
rlabel metal1 14766 12886 14766 12886 0 _093_
rlabel metal1 14582 12954 14582 12954 0 _094_
rlabel metal2 13294 14892 13294 14892 0 _095_
rlabel metal2 14122 11016 14122 11016 0 _096_
rlabel metal2 13938 10438 13938 10438 0 _097_
rlabel metal2 14214 10846 14214 10846 0 _098_
rlabel metal1 13708 13906 13708 13906 0 _099_
rlabel metal2 13570 4896 13570 4896 0 _100_
rlabel metal2 12742 7446 12742 7446 0 _101_
rlabel via1 12836 7378 12836 7378 0 _102_
rlabel metal1 13570 6970 13570 6970 0 _103_
rlabel metal1 13708 4590 13708 4590 0 _104_
rlabel metal2 11086 5542 11086 5542 0 _105_
rlabel metal1 10902 6664 10902 6664 0 _106_
rlabel metal1 11154 6766 11154 6766 0 _107_
rlabel metal1 11224 6426 11224 6426 0 _108_
rlabel metal2 10994 6154 10994 6154 0 _109_
rlabel metal1 14628 14450 14628 14450 0 _110_
rlabel metal1 14352 14858 14352 14858 0 _111_
rlabel metal2 12742 15249 12742 15249 0 _112_
rlabel via1 13386 12818 13386 12818 0 _113_
rlabel metal1 6348 14586 6348 14586 0 _114_
rlabel metal1 5888 12410 5888 12410 0 _115_
rlabel metal1 12650 10642 12650 10642 0 _116_
rlabel metal1 6233 12818 6233 12818 0 _117_
rlabel metal1 15226 13770 15226 13770 0 _118_
rlabel metal2 5842 13022 5842 13022 0 _119_
rlabel metal1 6256 12954 6256 12954 0 _120_
rlabel metal2 6210 9010 6210 9010 0 _121_
rlabel metal1 5934 10744 5934 10744 0 _122_
rlabel metal1 6233 10642 6233 10642 0 _123_
rlabel metal1 4968 10710 4968 10710 0 _124_
rlabel metal1 7912 9554 7912 9554 0 _125_
rlabel metal1 6072 4794 6072 4794 0 _126_
rlabel metal1 6348 5882 6348 5882 0 _127_
rlabel via1 6575 6290 6575 6290 0 _128_
rlabel metal1 5244 6358 5244 6358 0 _129_
rlabel metal2 6302 5882 6302 5882 0 _130_
rlabel metal1 10856 14994 10856 14994 0 _131_
rlabel metal1 10304 12274 10304 12274 0 _132_
rlabel via1 10623 13294 10623 13294 0 _133_
rlabel metal1 10810 13328 10810 13328 0 _134_
rlabel metal1 10488 13498 10488 13498 0 _135_
rlabel metal2 14766 14688 14766 14688 0 _136_
rlabel metal1 13662 12784 13662 12784 0 _137_
rlabel via1 13756 12818 13756 12818 0 _138_
rlabel metal2 13570 13464 13570 13464 0 _139_
rlabel metal1 14168 12954 14168 12954 0 _140_
rlabel metal2 14490 15606 14490 15606 0 _141_
rlabel metal1 13478 10608 13478 10608 0 _142_
rlabel via1 13572 10642 13572 10642 0 _143_
rlabel metal1 13708 10710 13708 10710 0 _144_
rlabel metal1 13892 14382 13892 14382 0 _145_
rlabel metal1 14628 4250 14628 4250 0 _146_
rlabel metal1 13248 7446 13248 7446 0 _147_
rlabel via1 13639 7378 13639 7378 0 _148_
rlabel metal1 13386 7344 13386 7344 0 _149_
rlabel metal1 14766 4624 14766 4624 0 _150_
rlabel metal1 11132 4794 11132 4794 0 _151_
rlabel metal2 11086 7038 11086 7038 0 _152_
rlabel via1 11180 6290 11180 6290 0 _153_
rlabel metal2 11362 6052 11362 6052 0 _154_
rlabel metal1 11500 5678 11500 5678 0 _155_
rlabel metal2 10810 9350 10810 9350 0 _156_
rlabel metal1 8050 16082 8050 16082 0 _157_
rlabel metal1 3726 15470 3726 15470 0 _158_
rlabel metal2 1794 9146 1794 9146 0 _159_
rlabel metal2 4554 5236 4554 5236 0 _160_
rlabel metal1 7452 16082 7452 16082 0 _161_
rlabel metal1 11408 14042 11408 14042 0 _162_
rlabel metal1 11546 16082 11546 16082 0 _163_
rlabel metal1 11592 4250 11592 4250 0 _164_
rlabel metal2 8326 4794 8326 4794 0 _165_
rlabel metal1 11086 9418 11086 9418 0 _166_
rlabel metal2 14674 2703 14674 2703 0 _167_
rlabel metal1 4922 16762 4922 16762 0 _168_
rlabel metal1 4140 8466 4140 8466 0 _169_
rlabel metal2 5842 3468 5842 3468 0 _170_
rlabel metal1 7958 17850 7958 17850 0 _171_
rlabel metal1 15318 17306 15318 17306 0 _172_
rlabel metal1 11684 17850 11684 17850 0 _173_
rlabel metal2 14122 3060 14122 3060 0 _174_
rlabel metal1 9476 3502 9476 3502 0 _175_
rlabel metal1 16054 15980 16054 15980 0 _176_
rlabel metal2 6026 17340 6026 17340 0 _177_
rlabel metal1 7636 8330 7636 8330 0 _178_
rlabel metal2 7866 2587 7866 2587 0 _179_
rlabel metal1 10304 17170 10304 17170 0 _180_
rlabel metal1 16376 14994 16376 14994 0 _181_
rlabel metal1 15410 16218 15410 16218 0 _182_
rlabel metal1 14720 3502 14720 3502 0 _183_
rlabel metal1 10166 3026 10166 3026 0 _184_
rlabel metal1 10672 8534 10672 8534 0 _185_
rlabel metal2 2668 12750 2668 12750 0 _186_
rlabel metal1 2070 12954 2070 12954 0 _187_
rlabel metal1 2116 10234 2116 10234 0 _188_
rlabel metal1 3312 4590 3312 4590 0 _189_
rlabel metal2 9338 14518 9338 14518 0 _190_
rlabel metal1 17434 13158 17434 13158 0 _191_
rlabel metal1 16284 10030 16284 10030 0 _192_
rlabel metal1 16698 6290 16698 6290 0 _193_
rlabel metal1 15226 4794 15226 4794 0 _194_
rlabel metal1 2484 11186 2484 11186 0 _195_
rlabel metal1 2254 14382 2254 14382 0 _196_
rlabel metal2 2070 11764 2070 11764 0 _197_
rlabel metal2 2898 6732 2898 6732 0 _198_
rlabel metal1 7590 14042 7590 14042 0 _199_
rlabel metal1 17066 14586 17066 14586 0 _200_
rlabel metal1 15594 11662 15594 11662 0 _201_
rlabel metal1 17296 8942 17296 8942 0 _202_
rlabel metal1 16468 5678 16468 5678 0 _203_
rlabel metal1 7912 8534 7912 8534 0 _204_
rlabel metal1 14766 10098 14766 10098 0 _205_
rlabel metal1 6854 12818 6854 12818 0 _206_
rlabel metal1 7360 10030 7360 10030 0 _207_
rlabel metal1 7912 6290 7912 6290 0 _208_
rlabel metal1 9844 10234 9844 10234 0 _209_
rlabel metal3 16468 12444 16468 12444 0 _210_
rlabel metal2 14858 10438 14858 10438 0 _211_
rlabel metal1 14996 8602 14996 8602 0 _212_
rlabel metal1 16192 6630 16192 6630 0 _213_
rlabel metal2 12144 12750 12144 12750 0 _214_
rlabel metal1 4232 12206 4232 12206 0 _215_
rlabel metal1 4232 11118 4232 11118 0 _216_
rlabel metal2 5474 7140 5474 7140 0 _217_
rlabel metal1 8740 11730 8740 11730 0 _218_
rlabel metal2 12650 13430 12650 13430 0 _219_
rlabel metal1 11592 10778 11592 10778 0 _220_
rlabel metal2 12006 9078 12006 9078 0 _221_
rlabel metal2 8970 6460 8970 6460 0 _222_
rlabel metal2 11454 9350 11454 9350 0 _223_
rlabel metal1 8234 17714 8234 17714 0 _224_
rlabel metal1 3496 16558 3496 16558 0 _225_
rlabel metal2 1886 8772 1886 8772 0 _226_
rlabel metal1 4508 3502 4508 3502 0 _227_
rlabel metal1 7176 17850 7176 17850 0 _228_
rlabel metal1 13892 17850 13892 17850 0 _229_
rlabel metal1 10948 17646 10948 17646 0 _230_
rlabel metal1 12880 3638 12880 3638 0 _231_
rlabel metal1 8970 3502 8970 3502 0 _232_
rlabel metal3 2131 17748 2131 17748 0 clk
rlabel metal1 13708 14314 13708 14314 0 clknet_0_clk
rlabel metal1 2622 5236 2622 5236 0 clknet_3_0__leaf_clk
rlabel metal1 8510 2482 8510 2482 0 clknet_3_1__leaf_clk
rlabel metal1 2622 17034 2622 17034 0 clknet_3_2__leaf_clk
rlabel metal1 8050 10676 8050 10676 0 clknet_3_3__leaf_clk
rlabel metal1 13202 6630 13202 6630 0 clknet_3_4__leaf_clk
rlabel metal1 14720 5134 14720 5134 0 clknet_3_5__leaf_clk
rlabel metal1 12857 18258 12857 18258 0 clknet_3_6__leaf_clk
rlabel metal2 15594 17136 15594 17136 0 clknet_3_7__leaf_clk
rlabel metal1 15180 5610 15180 5610 0 net1
rlabel metal1 4646 2550 4646 2550 0 net10
rlabel metal1 9384 13838 9384 13838 0 net11
rlabel metal2 14490 17408 14490 17408 0 net12
rlabel metal1 12052 17510 12052 17510 0 net13
rlabel metal1 14582 2516 14582 2516 0 net14
rlabel metal1 13524 2550 13524 2550 0 net15
rlabel metal1 11960 2482 11960 2482 0 net16
rlabel metal1 10856 2482 10856 2482 0 net17
rlabel metal1 8326 8908 8326 8908 0 net18
rlabel metal1 1702 15538 1702 15538 0 net19
rlabel metal1 14122 8432 14122 8432 0 net2
rlabel metal2 2070 9860 2070 9860 0 net20
rlabel metal1 6026 2414 6026 2414 0 net21
rlabel metal2 10534 16762 10534 16762 0 net22
rlabel metal1 15180 14586 15180 14586 0 net23
rlabel metal2 14122 16626 14122 16626 0 net24
rlabel metal1 17526 4692 17526 4692 0 net25
rlabel metal1 12880 2414 12880 2414 0 net26
rlabel metal1 1840 14382 1840 14382 0 net27
rlabel metal1 1702 9996 1702 9996 0 net28
rlabel metal1 6440 2414 6440 2414 0 net29
rlabel metal2 13294 13022 13294 13022 0 net3
rlabel metal1 9890 15130 9890 15130 0 net30
rlabel metal2 14674 13566 14674 13566 0 net31
rlabel metal1 16790 13838 16790 13838 0 net32
rlabel metal1 14398 4794 14398 4794 0 net33
rlabel metal1 12604 2414 12604 2414 0 net34
rlabel metal1 4462 8942 4462 8942 0 net35
rlabel metal1 4416 15470 4416 15470 0 net36
rlabel metal1 8418 16218 8418 16218 0 net37
rlabel metal1 12880 3434 12880 3434 0 net38
rlabel metal1 15824 15130 15824 15130 0 net39
rlabel metal1 14398 6834 14398 6834 0 net4
rlabel metal2 4646 11356 4646 11356 0 net40
rlabel metal2 2806 14620 2806 14620 0 net41
rlabel metal1 10856 16218 10856 16218 0 net42
rlabel metal2 2438 11594 2438 11594 0 net43
rlabel metal1 8878 5338 8878 5338 0 net44
rlabel metal1 12742 17646 12742 17646 0 net45
rlabel metal1 6992 4182 6992 4182 0 net46
rlabel metal1 3496 7378 3496 7378 0 net47
rlabel metal2 12742 4352 12742 4352 0 net48
rlabel metal1 11408 17646 11408 17646 0 net49
rlabel metal2 13478 8194 13478 8194 0 net5
rlabel metal1 5336 16490 5336 16490 0 net50
rlabel metal1 10672 3434 10672 3434 0 net51
rlabel metal1 16790 11730 16790 11730 0 net52
rlabel metal2 3818 8262 3818 8262 0 net53
rlabel metal2 8418 3706 8418 3706 0 net54
rlabel metal1 16422 14314 16422 14314 0 net55
rlabel metal1 4876 12138 4876 12138 0 net56
rlabel metal2 12098 10914 12098 10914 0 net57
rlabel metal1 9384 11730 9384 11730 0 net58
rlabel metal2 4922 3706 4922 3706 0 net59
rlabel metal2 1794 11934 1794 11934 0 net6
rlabel metal2 4186 17034 4186 17034 0 net60
rlabel metal1 9568 6766 9568 6766 0 net61
rlabel metal1 8694 17578 8694 17578 0 net62
rlabel metal2 12834 13022 12834 13022 0 net63
rlabel metal1 7268 8602 7268 8602 0 net64
rlabel metal1 5244 4590 5244 4590 0 net65
rlabel metal2 13202 8704 13202 8704 0 net66
rlabel metal1 7406 2618 7406 2618 0 net67
rlabel metal1 9844 17306 9844 17306 0 net68
rlabel metal2 12650 14688 12650 14688 0 net69
rlabel metal1 9292 8466 9292 8466 0 net7
rlabel metal1 2622 12954 2622 12954 0 net70
rlabel metal2 14582 17408 14582 17408 0 net71
rlabel metal1 15456 3434 15456 3434 0 net72
rlabel metal1 2484 9554 2484 9554 0 net73
rlabel metal1 14720 2346 14720 2346 0 net74
rlabel metal2 10994 3706 10994 3706 0 net75
rlabel metal1 16698 8942 16698 8942 0 net76
rlabel metal1 8142 14042 8142 14042 0 net77
rlabel metal1 7636 17646 7636 17646 0 net78
rlabel metal2 4186 10234 4186 10234 0 net79
rlabel metal1 2116 16626 2116 16626 0 net8
rlabel metal1 16468 16218 16468 16218 0 net80
rlabel metal1 14168 17578 14168 17578 0 net81
rlabel metal1 4416 5610 4416 5610 0 net82
rlabel metal2 17526 10438 17526 10438 0 net83
rlabel metal1 6440 17578 6440 17578 0 net84
rlabel metal2 8970 14110 8970 14110 0 net85
rlabel metal1 16652 4114 16652 4114 0 net86
rlabel metal1 15824 4114 15824 4114 0 net87
rlabel metal1 17066 13294 17066 13294 0 net88
rlabel metal1 5336 6290 5336 6290 0 net89
rlabel metal2 2714 9180 2714 9180 0 net9
rlabel metal1 15502 4590 15502 4590 0 net90
rlabel metal1 14674 9962 14674 9962 0 net91
rlabel metal1 7590 12308 7590 12308 0 net92
rlabel metal1 16284 12274 16284 12274 0 net93
rlabel metal1 7958 11050 7958 11050 0 net94
rlabel metal2 7314 7616 7314 7616 0 net95
rlabel metal2 15686 9010 15686 9010 0 net96
rlabel metal1 10626 9894 10626 9894 0 net97
rlabel metal2 15686 6528 15686 6528 0 net98
rlabel metal3 1096 15028 1096 15028 0 readData1[0]
rlabel metal3 1280 9588 1280 9588 0 readData1[1]
rlabel metal2 6486 1520 6486 1520 0 readData1[2]
rlabel metal1 9614 18394 9614 18394 0 readData1[3]
rlabel metal2 17710 15793 17710 15793 0 readData1[4]
rlabel metal2 12650 19839 12650 19839 0 readData1[5]
rlabel metal2 17710 5151 17710 5151 0 readData1[6]
rlabel metal2 11638 1656 11638 1656 0 readData1[7]
rlabel metal3 751 14348 751 14348 0 readData2[0]
rlabel metal1 1380 10234 1380 10234 0 readData2[1]
rlabel metal2 7130 1520 7130 1520 0 readData2[2]
rlabel metal1 10212 18938 10212 18938 0 readData2[3]
rlabel metal2 17710 15181 17710 15181 0 readData2[4]
rlabel metal2 16974 14195 16974 14195 0 readData2[5]
rlabel metal2 17618 4913 17618 4913 0 readData2[6]
rlabel metal2 10994 1520 10994 1520 0 readData2[7]
rlabel metal2 17802 5967 17802 5967 0 readReg1[0]
rlabel metal2 17802 7463 17802 7463 0 readReg1[1]
rlabel metal1 1288 12886 1288 12886 0 readReg1[2]
rlabel metal2 17802 6579 17802 6579 0 readReg2[0]
rlabel metal2 16974 8313 16974 8313 0 readReg2[1]
rlabel metal1 1426 12206 1426 12206 0 readReg2[2]
rlabel metal1 9246 3026 9246 3026 0 regWrite
rlabel metal1 7084 13294 7084 13294 0 registers\[0\]\[0\]
rlabel metal1 6992 11118 6992 11118 0 registers\[0\]\[1\]
rlabel metal1 7544 6970 7544 6970 0 registers\[0\]\[2\]
rlabel metal1 11224 12818 11224 12818 0 registers\[0\]\[3\]
rlabel metal1 15824 12614 15824 12614 0 registers\[0\]\[4\]
rlabel metal1 13570 10030 13570 10030 0 registers\[0\]\[5\]
rlabel metal2 16422 9316 16422 9316 0 registers\[0\]\[6\]
rlabel metal2 15042 6766 15042 6766 0 registers\[0\]\[7\]
rlabel metal1 5382 12954 5382 12954 0 registers\[1\]\[0\]
rlabel metal2 5382 11492 5382 11492 0 registers\[1\]\[1\]
rlabel via2 6210 6205 6210 6205 0 registers\[1\]\[2\]
rlabel metal1 9798 11662 9798 11662 0 registers\[1\]\[3\]
rlabel metal1 12742 13396 12742 13396 0 registers\[1\]\[4\]
rlabel metal2 12650 10710 12650 10710 0 registers\[1\]\[5\]
rlabel metal1 14076 9010 14076 9010 0 registers\[1\]\[6\]
rlabel metal2 10626 7072 10626 7072 0 registers\[1\]\[7\]
rlabel metal1 3542 14858 3542 14858 0 registers\[2\]\[0\]
rlabel metal2 3266 10880 3266 10880 0 registers\[2\]\[1\]
rlabel metal1 4232 6426 4232 6426 0 registers\[2\]\[2\]
rlabel metal1 8970 14892 8970 14892 0 registers\[2\]\[3\]
rlabel metal2 16422 14722 16422 14722 0 registers\[2\]\[4\]
rlabel metal1 15548 11118 15548 11118 0 registers\[2\]\[5\]
rlabel metal1 16376 8058 16376 8058 0 registers\[2\]\[6\]
rlabel metal1 12834 5678 12834 5678 0 registers\[2\]\[7\]
rlabel metal1 3312 13362 3312 13362 0 registers\[3\]\[0\]
rlabel metal1 4186 10642 4186 10642 0 registers\[3\]\[1\]
rlabel metal1 4094 6154 4094 6154 0 registers\[3\]\[2\]
rlabel viali 10362 14586 10362 14586 0 registers\[3\]\[3\]
rlabel metal1 16882 13974 16882 13974 0 registers\[3\]\[4\]
rlabel metal1 16468 10982 16468 10982 0 registers\[3\]\[5\]
rlabel metal1 17664 6630 17664 6630 0 registers\[3\]\[6\]
rlabel metal2 13294 6052 13294 6052 0 registers\[3\]\[7\]
rlabel metal1 4968 15470 4968 15470 0 registers\[4\]\[0\]
rlabel metal1 6854 9146 6854 9146 0 registers\[4\]\[1\]
rlabel via2 7314 4573 7314 4573 0 registers\[4\]\[2\]
rlabel metal1 10580 17850 10580 17850 0 registers\[4\]\[3\]
rlabel metal1 15824 15470 15824 15470 0 registers\[4\]\[4\]
rlabel metal1 17296 16558 17296 16558 0 registers\[4\]\[5\]
rlabel metal1 13064 4046 13064 4046 0 registers\[4\]\[6\]
rlabel metal1 9614 4658 9614 4658 0 registers\[4\]\[7\]
rlabel metal1 4784 15470 4784 15470 0 registers\[5\]\[0\]
rlabel metal1 4922 9452 4922 9452 0 registers\[5\]\[1\]
rlabel metal1 7452 4658 7452 4658 0 registers\[5\]\[2\]
rlabel metal2 9338 18564 9338 18564 0 registers\[5\]\[3\]
rlabel metal1 16330 17782 16330 17782 0 registers\[5\]\[4\]
rlabel metal2 13110 18564 13110 18564 0 registers\[5\]\[5\]
rlabel metal1 14352 2414 14352 2414 0 registers\[5\]\[6\]
rlabel metal1 10764 3570 10764 3570 0 registers\[5\]\[7\]
rlabel metal1 4876 16082 4876 16082 0 registers\[6\]\[0\]
rlabel metal2 2622 8908 2622 8908 0 registers\[6\]\[1\]
rlabel metal1 6440 5202 6440 5202 0 registers\[6\]\[2\]
rlabel metal1 9522 16660 9522 16660 0 registers\[6\]\[3\]
rlabel via1 13925 14994 13925 14994 0 registers\[6\]\[4\]
rlabel metal1 12800 16626 12800 16626 0 registers\[6\]\[5\]
rlabel metal1 13616 4658 13616 4658 0 registers\[6\]\[6\]
rlabel metal1 9522 5780 9522 5780 0 registers\[6\]\[7\]
rlabel metal2 4738 17476 4738 17476 0 registers\[7\]\[0\]
rlabel metal2 4370 8500 4370 8500 0 registers\[7\]\[1\]
rlabel metal1 5704 4046 5704 4046 0 registers\[7\]\[2\]
rlabel metal2 9522 15844 9522 15844 0 registers\[7\]\[3\]
rlabel metal2 15042 15232 15042 15232 0 registers\[7\]\[4\]
rlabel metal2 12650 18394 12650 18394 0 registers\[7\]\[5\]
rlabel metal2 13754 4658 13754 4658 0 registers\[7\]\[6\]
rlabel metal2 10166 4862 10166 4862 0 registers\[7\]\[7\]
rlabel metal3 751 16388 751 16388 0 writeData[0]
rlabel metal3 1096 10948 1096 10948 0 writeData[1]
rlabel metal2 3910 959 3910 959 0 writeData[2]
rlabel metal1 8878 18734 8878 18734 0 writeData[3]
rlabel metal2 17710 13107 17710 13107 0 writeData[4]
rlabel metal2 17710 10455 17710 10455 0 writeData[5]
rlabel via2 17710 3451 17710 3451 0 writeData[6]
rlabel metal2 12282 959 12282 959 0 writeData[7]
rlabel metal2 9706 1554 9706 1554 0 writeReg[0]
rlabel metal2 10350 1588 10350 1588 0 writeReg[1]
rlabel metal2 8418 1554 8418 1554 0 writeReg[2]
<< properties >>
string FIXED_BBOX 0 0 19269 21413
<< end >>
