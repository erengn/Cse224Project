module register_file (clk,
    regWrite,
    readData1,
    readData2,
    readReg1,
    readReg2,
    writeData,
    writeReg);
 input clk;
 input regWrite;
 output [7:0] readData1;
 output [7:0] readData2;
 input [2:0] readReg1;
 input [2:0] readReg2;
 input [7:0] writeData;
 input [2:0] writeReg;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire \registers[0][0] ;
 wire \registers[0][1] ;
 wire \registers[0][2] ;
 wire \registers[0][3] ;
 wire \registers[0][4] ;
 wire \registers[0][5] ;
 wire \registers[0][6] ;
 wire \registers[0][7] ;
 wire \registers[1][0] ;
 wire \registers[1][1] ;
 wire \registers[1][2] ;
 wire \registers[1][3] ;
 wire \registers[1][4] ;
 wire \registers[1][5] ;
 wire \registers[1][6] ;
 wire \registers[1][7] ;
 wire \registers[2][0] ;
 wire \registers[2][1] ;
 wire \registers[2][2] ;
 wire \registers[2][3] ;
 wire \registers[2][4] ;
 wire \registers[2][5] ;
 wire \registers[2][6] ;
 wire \registers[2][7] ;
 wire \registers[3][0] ;
 wire \registers[3][1] ;
 wire \registers[3][2] ;
 wire \registers[3][3] ;
 wire \registers[3][4] ;
 wire \registers[3][5] ;
 wire \registers[3][6] ;
 wire \registers[3][7] ;
 wire \registers[4][0] ;
 wire \registers[4][1] ;
 wire \registers[4][2] ;
 wire \registers[4][3] ;
 wire \registers[4][4] ;
 wire \registers[4][5] ;
 wire \registers[4][6] ;
 wire \registers[4][7] ;
 wire \registers[5][0] ;
 wire \registers[5][1] ;
 wire \registers[5][2] ;
 wire \registers[5][3] ;
 wire \registers[5][4] ;
 wire \registers[5][5] ;
 wire \registers[5][6] ;
 wire \registers[5][7] ;
 wire \registers[6][0] ;
 wire \registers[6][1] ;
 wire \registers[6][2] ;
 wire \registers[6][3] ;
 wire \registers[6][4] ;
 wire \registers[6][5] ;
 wire \registers[6][6] ;
 wire \registers[6][7] ;
 wire \registers[7][0] ;
 wire \registers[7][1] ;
 wire \registers[7][2] ;
 wire \registers[7][3] ;
 wire \registers[7][4] ;
 wire \registers[7][5] ;
 wire \registers[7][6] ;
 wire \registers[7][7] ;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;

 sky130_fd_sc_hd__inv_2 _233_ (.A(net6),
    .Y(_064_));
 sky130_fd_sc_hd__buf_4 _234_ (.A(net4),
    .X(_065_));
 sky130_fd_sc_hd__clkbuf_4 _235_ (.A(net5),
    .X(_066_));
 sky130_fd_sc_hd__clkbuf_4 _236_ (.A(_066_),
    .X(_067_));
 sky130_fd_sc_hd__mux4_1 _237_ (.A0(\registers[4][0] ),
    .A1(\registers[5][0] ),
    .A2(\registers[6][0] ),
    .A3(\registers[7][0] ),
    .S0(_065_),
    .S1(_067_),
    .X(_068_));
 sky130_fd_sc_hd__or2b_1 _238_ (.A(\registers[1][0] ),
    .B_N(_065_),
    .X(_069_));
 sky130_fd_sc_hd__buf_2 _239_ (.A(net4),
    .X(_070_));
 sky130_fd_sc_hd__o21ba_1 _240_ (.A1(\registers[0][0] ),
    .A2(_070_),
    .B1_N(_066_),
    .X(_071_));
 sky130_fd_sc_hd__clkbuf_4 _241_ (.A(net4),
    .X(_072_));
 sky130_fd_sc_hd__mux2_1 _242_ (.A0(\registers[2][0] ),
    .A1(\registers[3][0] ),
    .S(_072_),
    .X(_073_));
 sky130_fd_sc_hd__a221o_1 _243_ (.A1(_069_),
    .A2(_071_),
    .B1(_073_),
    .B2(_067_),
    .C1(net6),
    .X(_074_));
 sky130_fd_sc_hd__o21a_1 _244_ (.A1(_064_),
    .A2(_068_),
    .B1(_074_),
    .X(net27));
 sky130_fd_sc_hd__mux4_1 _245_ (.A0(\registers[4][1] ),
    .A1(\registers[5][1] ),
    .A2(\registers[6][1] ),
    .A3(\registers[7][1] ),
    .S0(_065_),
    .S1(_067_),
    .X(_075_));
 sky130_fd_sc_hd__or2b_1 _246_ (.A(\registers[1][1] ),
    .B_N(_065_),
    .X(_076_));
 sky130_fd_sc_hd__o21ba_1 _247_ (.A1(_070_),
    .A2(\registers[0][1] ),
    .B1_N(_066_),
    .X(_077_));
 sky130_fd_sc_hd__mux2_1 _248_ (.A0(\registers[2][1] ),
    .A1(\registers[3][1] ),
    .S(_072_),
    .X(_078_));
 sky130_fd_sc_hd__a221o_1 _249_ (.A1(_076_),
    .A2(_077_),
    .B1(_078_),
    .B2(_067_),
    .C1(net6),
    .X(_079_));
 sky130_fd_sc_hd__o21a_1 _250_ (.A1(_064_),
    .A2(_075_),
    .B1(_079_),
    .X(net28));
 sky130_fd_sc_hd__mux4_1 _251_ (.A0(\registers[4][2] ),
    .A1(\registers[5][2] ),
    .A2(\registers[6][2] ),
    .A3(\registers[7][2] ),
    .S0(_065_),
    .S1(_066_),
    .X(_080_));
 sky130_fd_sc_hd__or2b_1 _252_ (.A(\registers[1][2] ),
    .B_N(_070_),
    .X(_081_));
 sky130_fd_sc_hd__o21ba_1 _253_ (.A1(_070_),
    .A2(\registers[0][2] ),
    .B1_N(_066_),
    .X(_082_));
 sky130_fd_sc_hd__mux2_1 _254_ (.A0(\registers[2][2] ),
    .A1(\registers[3][2] ),
    .S(_072_),
    .X(_083_));
 sky130_fd_sc_hd__a221o_1 _255_ (.A1(_081_),
    .A2(_082_),
    .B1(_083_),
    .B2(_067_),
    .C1(net6),
    .X(_084_));
 sky130_fd_sc_hd__o21a_1 _256_ (.A1(_064_),
    .A2(_080_),
    .B1(_084_),
    .X(net29));
 sky130_fd_sc_hd__mux4_1 _257_ (.A0(\registers[4][3] ),
    .A1(\registers[5][3] ),
    .A2(\registers[6][3] ),
    .A3(\registers[7][3] ),
    .S0(_065_),
    .S1(_066_),
    .X(_085_));
 sky130_fd_sc_hd__or2b_1 _258_ (.A(\registers[1][3] ),
    .B_N(_070_),
    .X(_086_));
 sky130_fd_sc_hd__o21ba_1 _259_ (.A1(_070_),
    .A2(\registers[0][3] ),
    .B1_N(net5),
    .X(_087_));
 sky130_fd_sc_hd__mux2_1 _260_ (.A0(\registers[2][3] ),
    .A1(\registers[3][3] ),
    .S(_072_),
    .X(_088_));
 sky130_fd_sc_hd__a221o_1 _261_ (.A1(_086_),
    .A2(_087_),
    .B1(_088_),
    .B2(_067_),
    .C1(net6),
    .X(_089_));
 sky130_fd_sc_hd__o21a_1 _262_ (.A1(_064_),
    .A2(_085_),
    .B1(_089_),
    .X(net30));
 sky130_fd_sc_hd__mux4_1 _263_ (.A0(\registers[4][4] ),
    .A1(\registers[5][4] ),
    .A2(\registers[6][4] ),
    .A3(\registers[7][4] ),
    .S0(_065_),
    .S1(_066_),
    .X(_090_));
 sky130_fd_sc_hd__or2b_1 _264_ (.A(\registers[1][4] ),
    .B_N(_070_),
    .X(_091_));
 sky130_fd_sc_hd__o21ba_1 _265_ (.A1(_072_),
    .A2(\registers[0][4] ),
    .B1_N(net5),
    .X(_092_));
 sky130_fd_sc_hd__mux2_1 _266_ (.A0(\registers[2][4] ),
    .A1(\registers[3][4] ),
    .S(_072_),
    .X(_093_));
 sky130_fd_sc_hd__a221o_1 _267_ (.A1(_091_),
    .A2(_092_),
    .B1(_093_),
    .B2(_067_),
    .C1(net6),
    .X(_094_));
 sky130_fd_sc_hd__o21a_1 _268_ (.A1(_064_),
    .A2(_090_),
    .B1(_094_),
    .X(net31));
 sky130_fd_sc_hd__mux4_1 _269_ (.A0(\registers[4][5] ),
    .A1(\registers[5][5] ),
    .A2(\registers[6][5] ),
    .A3(\registers[7][5] ),
    .S0(_065_),
    .S1(_066_),
    .X(_095_));
 sky130_fd_sc_hd__or2b_1 _270_ (.A(\registers[1][5] ),
    .B_N(_070_),
    .X(_096_));
 sky130_fd_sc_hd__o21ba_1 _271_ (.A1(_072_),
    .A2(\registers[0][5] ),
    .B1_N(net5),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _272_ (.A0(\registers[2][5] ),
    .A1(\registers[3][5] ),
    .S(_072_),
    .X(_098_));
 sky130_fd_sc_hd__a221o_1 _273_ (.A1(_096_),
    .A2(_097_),
    .B1(_098_),
    .B2(_067_),
    .C1(net6),
    .X(_099_));
 sky130_fd_sc_hd__o21a_1 _274_ (.A1(_064_),
    .A2(_095_),
    .B1(_099_),
    .X(net32));
 sky130_fd_sc_hd__mux4_1 _275_ (.A0(\registers[4][6] ),
    .A1(\registers[5][6] ),
    .A2(\registers[6][6] ),
    .A3(\registers[7][6] ),
    .S0(_065_),
    .S1(_066_),
    .X(_100_));
 sky130_fd_sc_hd__or2b_1 _276_ (.A(\registers[1][6] ),
    .B_N(_070_),
    .X(_101_));
 sky130_fd_sc_hd__o21ba_1 _277_ (.A1(_072_),
    .A2(\registers[0][6] ),
    .B1_N(net5),
    .X(_102_));
 sky130_fd_sc_hd__mux2_1 _278_ (.A0(\registers[2][6] ),
    .A1(\registers[3][6] ),
    .S(net4),
    .X(_103_));
 sky130_fd_sc_hd__a221o_1 _279_ (.A1(_101_),
    .A2(_102_),
    .B1(_103_),
    .B2(_067_),
    .C1(net6),
    .X(_104_));
 sky130_fd_sc_hd__o21a_1 _280_ (.A1(_064_),
    .A2(_100_),
    .B1(_104_),
    .X(net33));
 sky130_fd_sc_hd__mux4_1 _281_ (.A0(\registers[4][7] ),
    .A1(\registers[5][7] ),
    .A2(\registers[6][7] ),
    .A3(\registers[7][7] ),
    .S0(_065_),
    .S1(_066_),
    .X(_105_));
 sky130_fd_sc_hd__or2b_1 _282_ (.A(\registers[1][7] ),
    .B_N(_070_),
    .X(_106_));
 sky130_fd_sc_hd__o21ba_1 _283_ (.A1(_072_),
    .A2(\registers[0][7] ),
    .B1_N(net5),
    .X(_107_));
 sky130_fd_sc_hd__mux2_1 _284_ (.A0(\registers[2][7] ),
    .A1(\registers[3][7] ),
    .S(net4),
    .X(_108_));
 sky130_fd_sc_hd__a221o_1 _285_ (.A1(_106_),
    .A2(_107_),
    .B1(_108_),
    .B2(_067_),
    .C1(net6),
    .X(_109_));
 sky130_fd_sc_hd__o21a_1 _286_ (.A1(_064_),
    .A2(_105_),
    .B1(_109_),
    .X(net34));
 sky130_fd_sc_hd__inv_2 _287_ (.A(net3),
    .Y(_110_));
 sky130_fd_sc_hd__buf_4 _288_ (.A(net1),
    .X(_111_));
 sky130_fd_sc_hd__clkbuf_4 _289_ (.A(net2),
    .X(_112_));
 sky130_fd_sc_hd__clkbuf_4 _290_ (.A(_112_),
    .X(_113_));
 sky130_fd_sc_hd__mux4_1 _291_ (.A0(\registers[4][0] ),
    .A1(\registers[5][0] ),
    .A2(\registers[6][0] ),
    .A3(\registers[7][0] ),
    .S0(_111_),
    .S1(_113_),
    .X(_114_));
 sky130_fd_sc_hd__or2b_1 _292_ (.A(\registers[1][0] ),
    .B_N(_111_),
    .X(_115_));
 sky130_fd_sc_hd__buf_2 _293_ (.A(net1),
    .X(_116_));
 sky130_fd_sc_hd__o21ba_1 _294_ (.A1(\registers[0][0] ),
    .A2(_116_),
    .B1_N(_112_),
    .X(_117_));
 sky130_fd_sc_hd__clkbuf_4 _295_ (.A(net1),
    .X(_118_));
 sky130_fd_sc_hd__mux2_1 _296_ (.A0(\registers[2][0] ),
    .A1(\registers[3][0] ),
    .S(_118_),
    .X(_119_));
 sky130_fd_sc_hd__a221o_1 _297_ (.A1(_115_),
    .A2(_117_),
    .B1(_119_),
    .B2(_113_),
    .C1(net3),
    .X(_120_));
 sky130_fd_sc_hd__o21a_1 _298_ (.A1(_110_),
    .A2(_114_),
    .B1(_120_),
    .X(net19));
 sky130_fd_sc_hd__mux4_1 _299_ (.A0(\registers[4][1] ),
    .A1(\registers[5][1] ),
    .A2(\registers[6][1] ),
    .A3(\registers[7][1] ),
    .S0(_111_),
    .S1(_113_),
    .X(_121_));
 sky130_fd_sc_hd__or2b_1 _300_ (.A(\registers[1][1] ),
    .B_N(_111_),
    .X(_122_));
 sky130_fd_sc_hd__o21ba_1 _301_ (.A1(\registers[0][1] ),
    .A2(_116_),
    .B1_N(_112_),
    .X(_123_));
 sky130_fd_sc_hd__mux2_1 _302_ (.A0(\registers[2][1] ),
    .A1(\registers[3][1] ),
    .S(_118_),
    .X(_124_));
 sky130_fd_sc_hd__a221o_1 _303_ (.A1(_122_),
    .A2(_123_),
    .B1(_124_),
    .B2(_113_),
    .C1(net3),
    .X(_125_));
 sky130_fd_sc_hd__o21a_1 _304_ (.A1(_110_),
    .A2(_121_),
    .B1(_125_),
    .X(net20));
 sky130_fd_sc_hd__mux4_1 _305_ (.A0(\registers[4][2] ),
    .A1(\registers[5][2] ),
    .A2(\registers[6][2] ),
    .A3(\registers[7][2] ),
    .S0(_111_),
    .S1(_112_),
    .X(_126_));
 sky130_fd_sc_hd__or2b_1 _306_ (.A(\registers[1][2] ),
    .B_N(_116_),
    .X(_127_));
 sky130_fd_sc_hd__o21ba_1 _307_ (.A1(\registers[0][2] ),
    .A2(_116_),
    .B1_N(_112_),
    .X(_128_));
 sky130_fd_sc_hd__mux2_1 _308_ (.A0(\registers[2][2] ),
    .A1(\registers[3][2] ),
    .S(_118_),
    .X(_129_));
 sky130_fd_sc_hd__a221o_1 _309_ (.A1(_127_),
    .A2(_128_),
    .B1(_129_),
    .B2(_113_),
    .C1(net3),
    .X(_130_));
 sky130_fd_sc_hd__o21a_1 _310_ (.A1(_110_),
    .A2(_126_),
    .B1(_130_),
    .X(net21));
 sky130_fd_sc_hd__mux4_1 _311_ (.A0(\registers[4][3] ),
    .A1(\registers[5][3] ),
    .A2(\registers[6][3] ),
    .A3(\registers[7][3] ),
    .S0(_111_),
    .S1(_112_),
    .X(_131_));
 sky130_fd_sc_hd__or2b_1 _312_ (.A(\registers[1][3] ),
    .B_N(_116_),
    .X(_132_));
 sky130_fd_sc_hd__o21ba_1 _313_ (.A1(\registers[0][3] ),
    .A2(_116_),
    .B1_N(net2),
    .X(_133_));
 sky130_fd_sc_hd__mux2_1 _314_ (.A0(\registers[2][3] ),
    .A1(\registers[3][3] ),
    .S(_118_),
    .X(_134_));
 sky130_fd_sc_hd__a221o_1 _315_ (.A1(_132_),
    .A2(_133_),
    .B1(_134_),
    .B2(_113_),
    .C1(net3),
    .X(_135_));
 sky130_fd_sc_hd__o21a_1 _316_ (.A1(_110_),
    .A2(_131_),
    .B1(_135_),
    .X(net22));
 sky130_fd_sc_hd__mux4_1 _317_ (.A0(\registers[4][4] ),
    .A1(\registers[5][4] ),
    .A2(\registers[6][4] ),
    .A3(\registers[7][4] ),
    .S0(_111_),
    .S1(_112_),
    .X(_136_));
 sky130_fd_sc_hd__or2b_1 _318_ (.A(\registers[1][4] ),
    .B_N(_116_),
    .X(_137_));
 sky130_fd_sc_hd__o21ba_1 _319_ (.A1(\registers[0][4] ),
    .A2(_118_),
    .B1_N(net2),
    .X(_138_));
 sky130_fd_sc_hd__mux2_1 _320_ (.A0(\registers[2][4] ),
    .A1(\registers[3][4] ),
    .S(_118_),
    .X(_139_));
 sky130_fd_sc_hd__a221o_1 _321_ (.A1(_137_),
    .A2(_138_),
    .B1(_139_),
    .B2(_113_),
    .C1(net3),
    .X(_140_));
 sky130_fd_sc_hd__o21a_1 _322_ (.A1(_110_),
    .A2(_136_),
    .B1(_140_),
    .X(net23));
 sky130_fd_sc_hd__mux4_1 _323_ (.A0(\registers[4][5] ),
    .A1(\registers[5][5] ),
    .A2(\registers[6][5] ),
    .A3(\registers[7][5] ),
    .S0(_111_),
    .S1(_112_),
    .X(_141_));
 sky130_fd_sc_hd__or2b_1 _324_ (.A(\registers[1][5] ),
    .B_N(_116_),
    .X(_142_));
 sky130_fd_sc_hd__o21ba_1 _325_ (.A1(\registers[0][5] ),
    .A2(_118_),
    .B1_N(net2),
    .X(_143_));
 sky130_fd_sc_hd__mux2_1 _326_ (.A0(\registers[2][5] ),
    .A1(\registers[3][5] ),
    .S(_118_),
    .X(_144_));
 sky130_fd_sc_hd__a221o_1 _327_ (.A1(_142_),
    .A2(_143_),
    .B1(_144_),
    .B2(_113_),
    .C1(net3),
    .X(_145_));
 sky130_fd_sc_hd__o21a_1 _328_ (.A1(_110_),
    .A2(_141_),
    .B1(_145_),
    .X(net24));
 sky130_fd_sc_hd__mux4_1 _329_ (.A0(\registers[4][6] ),
    .A1(\registers[5][6] ),
    .A2(\registers[6][6] ),
    .A3(\registers[7][6] ),
    .S0(_111_),
    .S1(_112_),
    .X(_146_));
 sky130_fd_sc_hd__or2b_1 _330_ (.A(\registers[1][6] ),
    .B_N(_116_),
    .X(_147_));
 sky130_fd_sc_hd__o21ba_1 _331_ (.A1(\registers[0][6] ),
    .A2(_118_),
    .B1_N(net2),
    .X(_148_));
 sky130_fd_sc_hd__mux2_1 _332_ (.A0(\registers[2][6] ),
    .A1(\registers[3][6] ),
    .S(net1),
    .X(_149_));
 sky130_fd_sc_hd__a221o_1 _333_ (.A1(_147_),
    .A2(_148_),
    .B1(_149_),
    .B2(_113_),
    .C1(net3),
    .X(_150_));
 sky130_fd_sc_hd__o21a_1 _334_ (.A1(_110_),
    .A2(_146_),
    .B1(_150_),
    .X(net25));
 sky130_fd_sc_hd__mux4_1 _335_ (.A0(\registers[4][7] ),
    .A1(\registers[5][7] ),
    .A2(\registers[6][7] ),
    .A3(\registers[7][7] ),
    .S0(_111_),
    .S1(_112_),
    .X(_151_));
 sky130_fd_sc_hd__or2b_1 _336_ (.A(\registers[1][7] ),
    .B_N(_116_),
    .X(_152_));
 sky130_fd_sc_hd__o21ba_1 _337_ (.A1(\registers[0][7] ),
    .A2(_118_),
    .B1_N(net2),
    .X(_153_));
 sky130_fd_sc_hd__mux2_1 _338_ (.A0(\registers[2][7] ),
    .A1(\registers[3][7] ),
    .S(net1),
    .X(_154_));
 sky130_fd_sc_hd__a221o_1 _339_ (.A1(_152_),
    .A2(_153_),
    .B1(_154_),
    .B2(_113_),
    .C1(net3),
    .X(_155_));
 sky130_fd_sc_hd__o21a_1 _340_ (.A1(_110_),
    .A2(_151_),
    .B1(_155_),
    .X(net26));
 sky130_fd_sc_hd__and4b_1 _341_ (.A_N(net16),
    .B(net7),
    .C(net18),
    .D(net17),
    .X(_156_));
 sky130_fd_sc_hd__clkbuf_4 _342_ (.A(_156_),
    .X(_157_));
 sky130_fd_sc_hd__mux2_1 _343_ (.A0(\registers[6][0] ),
    .A1(net8),
    .S(_157_),
    .X(_158_));
 sky130_fd_sc_hd__clkbuf_1 _344_ (.A(_158_),
    .X(_000_));
 sky130_fd_sc_hd__mux2_1 _345_ (.A0(\registers[6][1] ),
    .A1(net9),
    .S(_157_),
    .X(_159_));
 sky130_fd_sc_hd__clkbuf_1 _346_ (.A(_159_),
    .X(_001_));
 sky130_fd_sc_hd__mux2_1 _347_ (.A0(\registers[6][2] ),
    .A1(net10),
    .S(_157_),
    .X(_160_));
 sky130_fd_sc_hd__clkbuf_1 _348_ (.A(_160_),
    .X(_002_));
 sky130_fd_sc_hd__mux2_1 _349_ (.A0(\registers[6][3] ),
    .A1(net11),
    .S(_157_),
    .X(_161_));
 sky130_fd_sc_hd__clkbuf_1 _350_ (.A(_161_),
    .X(_003_));
 sky130_fd_sc_hd__mux2_1 _351_ (.A0(\registers[6][4] ),
    .A1(net12),
    .S(_157_),
    .X(_162_));
 sky130_fd_sc_hd__clkbuf_1 _352_ (.A(_162_),
    .X(_004_));
 sky130_fd_sc_hd__mux2_1 _353_ (.A0(\registers[6][5] ),
    .A1(net13),
    .S(_157_),
    .X(_163_));
 sky130_fd_sc_hd__clkbuf_1 _354_ (.A(_163_),
    .X(_005_));
 sky130_fd_sc_hd__mux2_1 _355_ (.A0(\registers[6][6] ),
    .A1(net14),
    .S(_157_),
    .X(_164_));
 sky130_fd_sc_hd__clkbuf_1 _356_ (.A(_164_),
    .X(_006_));
 sky130_fd_sc_hd__mux2_1 _357_ (.A0(\registers[6][7] ),
    .A1(net15),
    .S(_157_),
    .X(_165_));
 sky130_fd_sc_hd__clkbuf_1 _358_ (.A(_165_),
    .X(_007_));
 sky130_fd_sc_hd__and4b_1 _359_ (.A_N(net17),
    .B(net16),
    .C(net7),
    .D(net18),
    .X(_166_));
 sky130_fd_sc_hd__clkbuf_4 _360_ (.A(_166_),
    .X(_167_));
 sky130_fd_sc_hd__mux2_1 _361_ (.A0(\registers[5][0] ),
    .A1(net8),
    .S(_167_),
    .X(_168_));
 sky130_fd_sc_hd__clkbuf_1 _362_ (.A(_168_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _363_ (.A0(\registers[5][1] ),
    .A1(net9),
    .S(_167_),
    .X(_169_));
 sky130_fd_sc_hd__clkbuf_1 _364_ (.A(_169_),
    .X(_009_));
 sky130_fd_sc_hd__mux2_1 _365_ (.A0(\registers[5][2] ),
    .A1(net10),
    .S(_167_),
    .X(_170_));
 sky130_fd_sc_hd__clkbuf_1 _366_ (.A(_170_),
    .X(_010_));
 sky130_fd_sc_hd__mux2_1 _367_ (.A0(\registers[5][3] ),
    .A1(net11),
    .S(_167_),
    .X(_171_));
 sky130_fd_sc_hd__clkbuf_1 _368_ (.A(_171_),
    .X(_011_));
 sky130_fd_sc_hd__mux2_1 _369_ (.A0(\registers[5][4] ),
    .A1(net12),
    .S(_167_),
    .X(_172_));
 sky130_fd_sc_hd__clkbuf_1 _370_ (.A(_172_),
    .X(_012_));
 sky130_fd_sc_hd__mux2_1 _371_ (.A0(\registers[5][5] ),
    .A1(net13),
    .S(_167_),
    .X(_173_));
 sky130_fd_sc_hd__clkbuf_1 _372_ (.A(_173_),
    .X(_013_));
 sky130_fd_sc_hd__mux2_1 _373_ (.A0(\registers[5][6] ),
    .A1(net14),
    .S(_167_),
    .X(_174_));
 sky130_fd_sc_hd__clkbuf_1 _374_ (.A(_174_),
    .X(_014_));
 sky130_fd_sc_hd__mux2_1 _375_ (.A0(\registers[5][7] ),
    .A1(net15),
    .S(_167_),
    .X(_175_));
 sky130_fd_sc_hd__clkbuf_1 _376_ (.A(_175_),
    .X(_015_));
 sky130_fd_sc_hd__and4bb_4 _377_ (.A_N(net17),
    .B_N(net16),
    .C(net7),
    .D(net18),
    .X(_176_));
 sky130_fd_sc_hd__mux2_1 _378_ (.A0(\registers[4][0] ),
    .A1(net8),
    .S(_176_),
    .X(_177_));
 sky130_fd_sc_hd__clkbuf_1 _379_ (.A(_177_),
    .X(_016_));
 sky130_fd_sc_hd__mux2_1 _380_ (.A0(\registers[4][1] ),
    .A1(net9),
    .S(_176_),
    .X(_178_));
 sky130_fd_sc_hd__clkbuf_1 _381_ (.A(_178_),
    .X(_017_));
 sky130_fd_sc_hd__mux2_1 _382_ (.A0(\registers[4][2] ),
    .A1(net10),
    .S(_176_),
    .X(_179_));
 sky130_fd_sc_hd__clkbuf_1 _383_ (.A(_179_),
    .X(_018_));
 sky130_fd_sc_hd__mux2_1 _384_ (.A0(\registers[4][3] ),
    .A1(net11),
    .S(_176_),
    .X(_180_));
 sky130_fd_sc_hd__clkbuf_1 _385_ (.A(_180_),
    .X(_019_));
 sky130_fd_sc_hd__mux2_1 _386_ (.A0(\registers[4][4] ),
    .A1(net12),
    .S(_176_),
    .X(_181_));
 sky130_fd_sc_hd__clkbuf_1 _387_ (.A(_181_),
    .X(_020_));
 sky130_fd_sc_hd__mux2_1 _388_ (.A0(\registers[4][5] ),
    .A1(net13),
    .S(_176_),
    .X(_182_));
 sky130_fd_sc_hd__clkbuf_1 _389_ (.A(_182_),
    .X(_021_));
 sky130_fd_sc_hd__mux2_1 _390_ (.A0(\registers[4][6] ),
    .A1(net14),
    .S(_176_),
    .X(_183_));
 sky130_fd_sc_hd__clkbuf_1 _391_ (.A(_183_),
    .X(_022_));
 sky130_fd_sc_hd__mux2_1 _392_ (.A0(\registers[4][7] ),
    .A1(net15),
    .S(_176_),
    .X(_184_));
 sky130_fd_sc_hd__clkbuf_1 _393_ (.A(_184_),
    .X(_023_));
 sky130_fd_sc_hd__and4b_1 _394_ (.A_N(net18),
    .B(net17),
    .C(net16),
    .D(net7),
    .X(_185_));
 sky130_fd_sc_hd__clkbuf_4 _395_ (.A(_185_),
    .X(_186_));
 sky130_fd_sc_hd__mux2_1 _396_ (.A0(\registers[3][0] ),
    .A1(net8),
    .S(_186_),
    .X(_187_));
 sky130_fd_sc_hd__clkbuf_1 _397_ (.A(_187_),
    .X(_024_));
 sky130_fd_sc_hd__mux2_1 _398_ (.A0(\registers[3][1] ),
    .A1(net9),
    .S(_186_),
    .X(_188_));
 sky130_fd_sc_hd__clkbuf_1 _399_ (.A(_188_),
    .X(_025_));
 sky130_fd_sc_hd__mux2_1 _400_ (.A0(\registers[3][2] ),
    .A1(net10),
    .S(_186_),
    .X(_189_));
 sky130_fd_sc_hd__clkbuf_1 _401_ (.A(_189_),
    .X(_026_));
 sky130_fd_sc_hd__mux2_1 _402_ (.A0(\registers[3][3] ),
    .A1(net11),
    .S(_186_),
    .X(_190_));
 sky130_fd_sc_hd__clkbuf_1 _403_ (.A(_190_),
    .X(_027_));
 sky130_fd_sc_hd__mux2_1 _404_ (.A0(\registers[3][4] ),
    .A1(net12),
    .S(_186_),
    .X(_191_));
 sky130_fd_sc_hd__clkbuf_1 _405_ (.A(_191_),
    .X(_028_));
 sky130_fd_sc_hd__mux2_1 _406_ (.A0(\registers[3][5] ),
    .A1(net13),
    .S(_186_),
    .X(_192_));
 sky130_fd_sc_hd__clkbuf_1 _407_ (.A(_192_),
    .X(_029_));
 sky130_fd_sc_hd__mux2_1 _408_ (.A0(\registers[3][6] ),
    .A1(net14),
    .S(_186_),
    .X(_193_));
 sky130_fd_sc_hd__clkbuf_1 _409_ (.A(_193_),
    .X(_030_));
 sky130_fd_sc_hd__mux2_1 _410_ (.A0(\registers[3][7] ),
    .A1(net15),
    .S(_186_),
    .X(_194_));
 sky130_fd_sc_hd__clkbuf_1 _411_ (.A(_194_),
    .X(_031_));
 sky130_fd_sc_hd__and4bb_4 _412_ (.A_N(net18),
    .B_N(net16),
    .C(net7),
    .D(net17),
    .X(_195_));
 sky130_fd_sc_hd__mux2_1 _413_ (.A0(\registers[2][0] ),
    .A1(net8),
    .S(_195_),
    .X(_196_));
 sky130_fd_sc_hd__clkbuf_1 _414_ (.A(_196_),
    .X(_032_));
 sky130_fd_sc_hd__mux2_1 _415_ (.A0(\registers[2][1] ),
    .A1(net9),
    .S(_195_),
    .X(_197_));
 sky130_fd_sc_hd__clkbuf_1 _416_ (.A(_197_),
    .X(_033_));
 sky130_fd_sc_hd__mux2_1 _417_ (.A0(\registers[2][2] ),
    .A1(net10),
    .S(_195_),
    .X(_198_));
 sky130_fd_sc_hd__clkbuf_1 _418_ (.A(_198_),
    .X(_034_));
 sky130_fd_sc_hd__mux2_1 _419_ (.A0(\registers[2][3] ),
    .A1(net11),
    .S(_195_),
    .X(_199_));
 sky130_fd_sc_hd__clkbuf_1 _420_ (.A(_199_),
    .X(_035_));
 sky130_fd_sc_hd__mux2_1 _421_ (.A0(\registers[2][4] ),
    .A1(net12),
    .S(_195_),
    .X(_200_));
 sky130_fd_sc_hd__clkbuf_1 _422_ (.A(_200_),
    .X(_036_));
 sky130_fd_sc_hd__mux2_1 _423_ (.A0(\registers[2][5] ),
    .A1(net13),
    .S(_195_),
    .X(_201_));
 sky130_fd_sc_hd__clkbuf_1 _424_ (.A(_201_),
    .X(_037_));
 sky130_fd_sc_hd__mux2_1 _425_ (.A0(\registers[2][6] ),
    .A1(net14),
    .S(_195_),
    .X(_202_));
 sky130_fd_sc_hd__clkbuf_1 _426_ (.A(_202_),
    .X(_038_));
 sky130_fd_sc_hd__mux2_1 _427_ (.A0(\registers[2][7] ),
    .A1(net15),
    .S(_195_),
    .X(_203_));
 sky130_fd_sc_hd__clkbuf_1 _428_ (.A(_203_),
    .X(_039_));
 sky130_fd_sc_hd__or4b_1 _429_ (.A(net18),
    .B(net17),
    .C(net16),
    .D_N(net7),
    .X(_204_));
 sky130_fd_sc_hd__clkbuf_4 _430_ (.A(_204_),
    .X(_205_));
 sky130_fd_sc_hd__mux2_1 _431_ (.A0(net8),
    .A1(\registers[0][0] ),
    .S(_205_),
    .X(_206_));
 sky130_fd_sc_hd__clkbuf_1 _432_ (.A(_206_),
    .X(_040_));
 sky130_fd_sc_hd__mux2_1 _433_ (.A0(net9),
    .A1(\registers[0][1] ),
    .S(_205_),
    .X(_207_));
 sky130_fd_sc_hd__clkbuf_1 _434_ (.A(_207_),
    .X(_041_));
 sky130_fd_sc_hd__mux2_1 _435_ (.A0(net10),
    .A1(\registers[0][2] ),
    .S(_205_),
    .X(_208_));
 sky130_fd_sc_hd__clkbuf_1 _436_ (.A(_208_),
    .X(_042_));
 sky130_fd_sc_hd__mux2_1 _437_ (.A0(net11),
    .A1(\registers[0][3] ),
    .S(_205_),
    .X(_209_));
 sky130_fd_sc_hd__clkbuf_1 _438_ (.A(_209_),
    .X(_043_));
 sky130_fd_sc_hd__mux2_1 _439_ (.A0(net12),
    .A1(\registers[0][4] ),
    .S(_205_),
    .X(_210_));
 sky130_fd_sc_hd__clkbuf_1 _440_ (.A(_210_),
    .X(_044_));
 sky130_fd_sc_hd__mux2_1 _441_ (.A0(net13),
    .A1(\registers[0][5] ),
    .S(_205_),
    .X(_211_));
 sky130_fd_sc_hd__clkbuf_1 _442_ (.A(_211_),
    .X(_045_));
 sky130_fd_sc_hd__mux2_1 _443_ (.A0(net14),
    .A1(\registers[0][6] ),
    .S(_205_),
    .X(_212_));
 sky130_fd_sc_hd__clkbuf_1 _444_ (.A(_212_),
    .X(_046_));
 sky130_fd_sc_hd__mux2_1 _445_ (.A0(net15),
    .A1(\registers[0][7] ),
    .S(_205_),
    .X(_213_));
 sky130_fd_sc_hd__clkbuf_1 _446_ (.A(_213_),
    .X(_047_));
 sky130_fd_sc_hd__and4bb_4 _447_ (.A_N(net18),
    .B_N(net17),
    .C(net16),
    .D(net7),
    .X(_214_));
 sky130_fd_sc_hd__mux2_1 _448_ (.A0(\registers[1][0] ),
    .A1(net8),
    .S(_214_),
    .X(_215_));
 sky130_fd_sc_hd__clkbuf_1 _449_ (.A(_215_),
    .X(_048_));
 sky130_fd_sc_hd__mux2_1 _450_ (.A0(\registers[1][1] ),
    .A1(net9),
    .S(_214_),
    .X(_216_));
 sky130_fd_sc_hd__clkbuf_1 _451_ (.A(_216_),
    .X(_049_));
 sky130_fd_sc_hd__mux2_1 _452_ (.A0(\registers[1][2] ),
    .A1(net10),
    .S(_214_),
    .X(_217_));
 sky130_fd_sc_hd__clkbuf_1 _453_ (.A(_217_),
    .X(_050_));
 sky130_fd_sc_hd__mux2_1 _454_ (.A0(\registers[1][3] ),
    .A1(net11),
    .S(_214_),
    .X(_218_));
 sky130_fd_sc_hd__clkbuf_1 _455_ (.A(_218_),
    .X(_051_));
 sky130_fd_sc_hd__mux2_1 _456_ (.A0(\registers[1][4] ),
    .A1(net12),
    .S(_214_),
    .X(_219_));
 sky130_fd_sc_hd__clkbuf_1 _457_ (.A(_219_),
    .X(_052_));
 sky130_fd_sc_hd__mux2_1 _458_ (.A0(\registers[1][5] ),
    .A1(net13),
    .S(_214_),
    .X(_220_));
 sky130_fd_sc_hd__clkbuf_1 _459_ (.A(_220_),
    .X(_053_));
 sky130_fd_sc_hd__mux2_1 _460_ (.A0(\registers[1][6] ),
    .A1(net14),
    .S(_214_),
    .X(_221_));
 sky130_fd_sc_hd__clkbuf_1 _461_ (.A(_221_),
    .X(_054_));
 sky130_fd_sc_hd__mux2_1 _462_ (.A0(\registers[1][7] ),
    .A1(net15),
    .S(_214_),
    .X(_222_));
 sky130_fd_sc_hd__clkbuf_1 _463_ (.A(_222_),
    .X(_055_));
 sky130_fd_sc_hd__and4_1 _464_ (.A(net18),
    .B(net17),
    .C(net16),
    .D(net7),
    .X(_223_));
 sky130_fd_sc_hd__clkbuf_4 _465_ (.A(_223_),
    .X(_224_));
 sky130_fd_sc_hd__mux2_1 _466_ (.A0(\registers[7][0] ),
    .A1(net8),
    .S(_224_),
    .X(_225_));
 sky130_fd_sc_hd__clkbuf_1 _467_ (.A(_225_),
    .X(_056_));
 sky130_fd_sc_hd__mux2_1 _468_ (.A0(\registers[7][1] ),
    .A1(net9),
    .S(_224_),
    .X(_226_));
 sky130_fd_sc_hd__clkbuf_1 _469_ (.A(_226_),
    .X(_057_));
 sky130_fd_sc_hd__mux2_1 _470_ (.A0(\registers[7][2] ),
    .A1(net10),
    .S(_224_),
    .X(_227_));
 sky130_fd_sc_hd__clkbuf_1 _471_ (.A(_227_),
    .X(_058_));
 sky130_fd_sc_hd__mux2_1 _472_ (.A0(\registers[7][3] ),
    .A1(net11),
    .S(_224_),
    .X(_228_));
 sky130_fd_sc_hd__clkbuf_1 _473_ (.A(_228_),
    .X(_059_));
 sky130_fd_sc_hd__mux2_1 _474_ (.A0(\registers[7][4] ),
    .A1(net12),
    .S(_224_),
    .X(_229_));
 sky130_fd_sc_hd__clkbuf_1 _475_ (.A(_229_),
    .X(_060_));
 sky130_fd_sc_hd__mux2_1 _476_ (.A0(\registers[7][5] ),
    .A1(net13),
    .S(_224_),
    .X(_230_));
 sky130_fd_sc_hd__clkbuf_1 _477_ (.A(_230_),
    .X(_061_));
 sky130_fd_sc_hd__mux2_1 _478_ (.A0(\registers[7][6] ),
    .A1(net14),
    .S(_224_),
    .X(_231_));
 sky130_fd_sc_hd__clkbuf_1 _479_ (.A(_231_),
    .X(_062_));
 sky130_fd_sc_hd__mux2_1 _480_ (.A0(\registers[7][7] ),
    .A1(net15),
    .S(_224_),
    .X(_232_));
 sky130_fd_sc_hd__clkbuf_1 _481_ (.A(_232_),
    .X(_063_));
 sky130_fd_sc_hd__dfxtp_1 _482_ (.CLK(clk),
    .D(_000_),
    .Q(\registers[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 _483_ (.CLK(clk),
    .D(_001_),
    .Q(\registers[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 _484_ (.CLK(clk),
    .D(_002_),
    .Q(\registers[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 _485_ (.CLK(clk),
    .D(_003_),
    .Q(\registers[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 _486_ (.CLK(clk),
    .D(_004_),
    .Q(\registers[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 _487_ (.CLK(clk),
    .D(_005_),
    .Q(\registers[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 _488_ (.CLK(clk),
    .D(_006_),
    .Q(\registers[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 _489_ (.CLK(clk),
    .D(_007_),
    .Q(\registers[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 _490_ (.CLK(clk),
    .D(_008_),
    .Q(\registers[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 _491_ (.CLK(clk),
    .D(_009_),
    .Q(\registers[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 _492_ (.CLK(clk),
    .D(_010_),
    .Q(\registers[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 _493_ (.CLK(clk),
    .D(_011_),
    .Q(\registers[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 _494_ (.CLK(clk),
    .D(_012_),
    .Q(\registers[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 _495_ (.CLK(clk),
    .D(_013_),
    .Q(\registers[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 _496_ (.CLK(clk),
    .D(_014_),
    .Q(\registers[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 _497_ (.CLK(clk),
    .D(_015_),
    .Q(\registers[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 _498_ (.CLK(clk),
    .D(_016_),
    .Q(\registers[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 _499_ (.CLK(clk),
    .D(_017_),
    .Q(\registers[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 _500_ (.CLK(clk),
    .D(_018_),
    .Q(\registers[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 _501_ (.CLK(clk),
    .D(_019_),
    .Q(\registers[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 _502_ (.CLK(clk),
    .D(_020_),
    .Q(\registers[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 _503_ (.CLK(clk),
    .D(_021_),
    .Q(\registers[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 _504_ (.CLK(clk),
    .D(_022_),
    .Q(\registers[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 _505_ (.CLK(clk),
    .D(_023_),
    .Q(\registers[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 _506_ (.CLK(clk),
    .D(_024_),
    .Q(\registers[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 _507_ (.CLK(clk),
    .D(_025_),
    .Q(\registers[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 _508_ (.CLK(clk),
    .D(_026_),
    .Q(\registers[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 _509_ (.CLK(clk),
    .D(_027_),
    .Q(\registers[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 _510_ (.CLK(clk),
    .D(_028_),
    .Q(\registers[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 _511_ (.CLK(clk),
    .D(_029_),
    .Q(\registers[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 _512_ (.CLK(clk),
    .D(_030_),
    .Q(\registers[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 _513_ (.CLK(clk),
    .D(_031_),
    .Q(\registers[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 _514_ (.CLK(clk),
    .D(_032_),
    .Q(\registers[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 _515_ (.CLK(clk),
    .D(_033_),
    .Q(\registers[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 _516_ (.CLK(clk),
    .D(_034_),
    .Q(\registers[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 _517_ (.CLK(clk),
    .D(_035_),
    .Q(\registers[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 _518_ (.CLK(clk),
    .D(_036_),
    .Q(\registers[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 _519_ (.CLK(clk),
    .D(_037_),
    .Q(\registers[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 _520_ (.CLK(clk),
    .D(_038_),
    .Q(\registers[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 _521_ (.CLK(clk),
    .D(_039_),
    .Q(\registers[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 _522_ (.CLK(clk),
    .D(_040_),
    .Q(\registers[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _523_ (.CLK(clk),
    .D(_041_),
    .Q(\registers[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _524_ (.CLK(clk),
    .D(_042_),
    .Q(\registers[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _525_ (.CLK(clk),
    .D(_043_),
    .Q(\registers[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _526_ (.CLK(clk),
    .D(_044_),
    .Q(\registers[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _527_ (.CLK(clk),
    .D(_045_),
    .Q(\registers[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _528_ (.CLK(clk),
    .D(_046_),
    .Q(\registers[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _529_ (.CLK(clk),
    .D(_047_),
    .Q(\registers[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _530_ (.CLK(clk),
    .D(_048_),
    .Q(\registers[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _531_ (.CLK(clk),
    .D(_049_),
    .Q(\registers[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _532_ (.CLK(clk),
    .D(_050_),
    .Q(\registers[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _533_ (.CLK(clk),
    .D(_051_),
    .Q(\registers[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _534_ (.CLK(clk),
    .D(_052_),
    .Q(\registers[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _535_ (.CLK(clk),
    .D(_053_),
    .Q(\registers[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _536_ (.CLK(clk),
    .D(_054_),
    .Q(\registers[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _537_ (.CLK(clk),
    .D(_055_),
    .Q(\registers[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _538_ (.CLK(clk),
    .D(_056_),
    .Q(\registers[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 _539_ (.CLK(clk),
    .D(_057_),
    .Q(\registers[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 _540_ (.CLK(clk),
    .D(_058_),
    .Q(\registers[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 _541_ (.CLK(clk),
    .D(_059_),
    .Q(\registers[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 _542_ (.CLK(clk),
    .D(_060_),
    .Q(\registers[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 _543_ (.CLK(clk),
    .D(_061_),
    .Q(\registers[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 _544_ (.CLK(clk),
    .D(_062_),
    .Q(\registers[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 _545_ (.CLK(clk),
    .D(_063_),
    .Q(\registers[7][7] ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_160 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(readReg1[0]),
    .X(net1));
 sky130_fd_sc_hd__dlymetal6s2s_1 input2 (.A(readReg1[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_4 input3 (.A(readReg1[2]),
    .X(net3));
 sky130_fd_sc_hd__dlymetal6s2s_1 input4 (.A(readReg2[0]),
    .X(net4));
 sky130_fd_sc_hd__dlymetal6s2s_1 input5 (.A(readReg2[1]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input6 (.A(readReg2[2]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(regWrite),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(writeData[0]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_2 input9 (.A(writeData[1]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 input10 (.A(writeData[2]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_2 input11 (.A(writeData[3]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 input12 (.A(writeData[4]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input13 (.A(writeData[5]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 input14 (.A(writeData[6]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 input15 (.A(writeData[7]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(writeReg[0]),
    .X(net16));
 sky130_fd_sc_hd__dlymetal6s2s_1 input17 (.A(writeReg[1]),
    .X(net17));
 sky130_fd_sc_hd__dlymetal6s2s_1 input18 (.A(writeReg[2]),
    .X(net18));
 sky130_fd_sc_hd__buf_2 output19 (.A(net19),
    .X(readData1[0]));
 sky130_fd_sc_hd__buf_2 output20 (.A(net20),
    .X(readData1[1]));
 sky130_fd_sc_hd__buf_2 output21 (.A(net21),
    .X(readData1[2]));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(readData1[3]));
 sky130_fd_sc_hd__buf_2 output23 (.A(net23),
    .X(readData1[4]));
 sky130_fd_sc_hd__clkbuf_4 output24 (.A(net24),
    .X(readData1[5]));
 sky130_fd_sc_hd__buf_2 output25 (.A(net25),
    .X(readData1[6]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(readData1[7]));
 sky130_fd_sc_hd__buf_2 output27 (.A(net27),
    .X(readData2[0]));
 sky130_fd_sc_hd__buf_2 output28 (.A(net28),
    .X(readData2[1]));
 sky130_fd_sc_hd__buf_2 output29 (.A(net29),
    .X(readData2[2]));
 sky130_fd_sc_hd__clkbuf_4 output30 (.A(net30),
    .X(readData2[3]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(readData2[4]));
 sky130_fd_sc_hd__buf_2 output32 (.A(net32),
    .X(readData2[5]));
 sky130_fd_sc_hd__buf_2 output33 (.A(net33),
    .X(readData2[6]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(readData2[7]));
endmodule
