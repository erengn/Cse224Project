# Temporary LEF after floorplan
